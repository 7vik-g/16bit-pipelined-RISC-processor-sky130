magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< locali >>
rect 70 282 136 316
rect 549 314 970 348
rect 70 174 136 208
rect 936 170 970 314
rect 1705 103 4122 137
<< metal1 >>
rect 246 -30 294 402
rect 670 -32 720 402
rect 1724 0 1752 395
rect 3372 0 3400 395
use sky130_fd_bd_sram__openram_dp_nand2_dec_1  sky130_fd_bd_sram__openram_dp_nand2_dec_0
timestamp 1666464484
transform 1 0 0 0 1 0
box 70 -56 888 476
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_dec_0  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_dec_0_0
timestamp 1666464484
transform 1 0 876 0 1 0
box 44 0 3264 490
<< labels >>
rlabel metal1 s 670 -32 720 402 4 vdd
port 1 nsew
rlabel metal1 s 3372 0 3400 395 4 vdd
port 1 nsew
rlabel metal1 s 246 -30 294 402 4 gnd
port 2 nsew
rlabel metal1 s 1724 0 1752 395 4 gnd
port 2 nsew
rlabel locali s 2913 120 2913 120 4 Z
port 3 nsew
rlabel locali s 103 299 103 299 4 A
port 4 nsew
rlabel locali s 103 191 103 191 4 B
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 4122 395
string GDS_END 151226
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 149738
<< end >>
