magic
tech sky130B
timestamp 1666464484
<< properties >>
string GDS_END 67584
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 67260
<< end >>
