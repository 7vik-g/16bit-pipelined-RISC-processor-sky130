magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< metal1 >>
rect 13910 1399 13916 1451
rect 13968 1399 13974 1451
rect 15158 1399 15164 1451
rect 15216 1399 15222 1451
rect 16406 1399 16412 1451
rect 16464 1399 16470 1451
rect 17654 1399 17660 1451
rect 17712 1399 17718 1451
rect 18902 1399 18908 1451
rect 18960 1399 18966 1451
rect 20150 1399 20156 1451
rect 20208 1399 20214 1451
rect 21398 1399 21404 1451
rect 21456 1399 21462 1451
rect 22646 1399 22652 1451
rect 22704 1399 22710 1451
rect 23894 1399 23900 1451
rect 23952 1399 23958 1451
rect 25142 1399 25148 1451
rect 25200 1399 25206 1451
rect 26390 1399 26396 1451
rect 26448 1399 26454 1451
rect 27638 1399 27644 1451
rect 27696 1399 27702 1451
rect 28886 1399 28892 1451
rect 28944 1399 28950 1451
rect 30134 1399 30140 1451
rect 30192 1399 30198 1451
rect 31382 1399 31388 1451
rect 31440 1399 31446 1451
rect 32630 1399 32636 1451
rect 32688 1399 32694 1451
rect 33878 1399 33884 1451
rect 33936 1399 33942 1451
rect 35126 1399 35132 1451
rect 35184 1399 35190 1451
rect 36374 1399 36380 1451
rect 36432 1399 36438 1451
rect 37622 1399 37628 1451
rect 37680 1399 37686 1451
rect 38870 1399 38876 1451
rect 38928 1399 38934 1451
rect 40118 1399 40124 1451
rect 40176 1399 40182 1451
rect 41366 1399 41372 1451
rect 41424 1399 41430 1451
rect 42614 1399 42620 1451
rect 42672 1399 42678 1451
rect 43862 1399 43868 1451
rect 43920 1399 43926 1451
rect 45110 1399 45116 1451
rect 45168 1399 45174 1451
rect 46358 1399 46364 1451
rect 46416 1399 46422 1451
rect 47606 1399 47612 1451
rect 47664 1399 47670 1451
rect 48854 1399 48860 1451
rect 48912 1399 48918 1451
rect 50102 1399 50108 1451
rect 50160 1399 50166 1451
rect 51350 1399 51356 1451
rect 51408 1399 51414 1451
rect 52598 1399 52604 1451
rect 52656 1399 52662 1451
<< via1 >>
rect 13916 1399 13968 1451
rect 15164 1399 15216 1451
rect 16412 1399 16464 1451
rect 17660 1399 17712 1451
rect 18908 1399 18960 1451
rect 20156 1399 20208 1451
rect 21404 1399 21456 1451
rect 22652 1399 22704 1451
rect 23900 1399 23952 1451
rect 25148 1399 25200 1451
rect 26396 1399 26448 1451
rect 27644 1399 27696 1451
rect 28892 1399 28944 1451
rect 30140 1399 30192 1451
rect 31388 1399 31440 1451
rect 32636 1399 32688 1451
rect 33884 1399 33936 1451
rect 35132 1399 35184 1451
rect 36380 1399 36432 1451
rect 37628 1399 37680 1451
rect 38876 1399 38928 1451
rect 40124 1399 40176 1451
rect 41372 1399 41424 1451
rect 42620 1399 42672 1451
rect 43868 1399 43920 1451
rect 45116 1399 45168 1451
rect 46364 1399 46416 1451
rect 47612 1399 47664 1451
rect 48860 1399 48912 1451
rect 50108 1399 50160 1451
rect 51356 1399 51408 1451
rect 52604 1399 52656 1451
<< metal2 >>
rect 13914 1453 13970 1462
rect 13914 1388 13970 1397
rect 15162 1453 15218 1462
rect 15162 1388 15218 1397
rect 16410 1453 16466 1462
rect 16410 1388 16466 1397
rect 17658 1453 17714 1462
rect 17658 1388 17714 1397
rect 18906 1453 18962 1462
rect 18906 1388 18962 1397
rect 20154 1453 20210 1462
rect 20154 1388 20210 1397
rect 21402 1453 21458 1462
rect 21402 1388 21458 1397
rect 22650 1453 22706 1462
rect 22650 1388 22706 1397
rect 23898 1453 23954 1462
rect 23898 1388 23954 1397
rect 25146 1453 25202 1462
rect 25146 1388 25202 1397
rect 26394 1453 26450 1462
rect 26394 1388 26450 1397
rect 27642 1453 27698 1462
rect 27642 1388 27698 1397
rect 28890 1453 28946 1462
rect 28890 1388 28946 1397
rect 30138 1453 30194 1462
rect 30138 1388 30194 1397
rect 31386 1453 31442 1462
rect 31386 1388 31442 1397
rect 32634 1453 32690 1462
rect 32634 1388 32690 1397
rect 33882 1453 33938 1462
rect 33882 1388 33938 1397
rect 35130 1453 35186 1462
rect 35130 1388 35186 1397
rect 36378 1453 36434 1462
rect 36378 1388 36434 1397
rect 37626 1453 37682 1462
rect 37626 1388 37682 1397
rect 38874 1453 38930 1462
rect 38874 1388 38930 1397
rect 40122 1453 40178 1462
rect 40122 1388 40178 1397
rect 41370 1453 41426 1462
rect 41370 1388 41426 1397
rect 42618 1453 42674 1462
rect 42618 1388 42674 1397
rect 43866 1453 43922 1462
rect 43866 1388 43922 1397
rect 45114 1453 45170 1462
rect 45114 1388 45170 1397
rect 46362 1453 46418 1462
rect 46362 1388 46418 1397
rect 47610 1453 47666 1462
rect 47610 1388 47666 1397
rect 48858 1453 48914 1462
rect 48858 1388 48914 1397
rect 50106 1453 50162 1462
rect 50106 1388 50162 1397
rect 51354 1453 51410 1462
rect 51354 1388 51410 1397
rect 52602 1453 52658 1462
rect 52602 1388 52658 1397
rect 13629 333 13685 342
rect 13629 268 13685 277
rect 23613 333 23669 342
rect 23613 268 23669 277
rect 33597 333 33653 342
rect 33597 268 33653 277
rect 43581 333 43637 342
rect 43581 268 43637 277
rect 3255 -3897 3311 -3888
rect 3255 -3962 3311 -3953
rect 4423 -3897 4479 -3888
rect 4423 -3962 4479 -3953
rect 5591 -3897 5647 -3888
rect 5591 -3962 5647 -3953
rect 6759 -3897 6815 -3888
rect 6759 -3962 6815 -3953
rect 7927 -3897 7983 -3888
rect 7927 -3962 7983 -3953
rect 9095 -3897 9151 -3888
rect 9095 -3962 9151 -3953
rect 10263 -3897 10319 -3888
rect 10263 -3962 10319 -3953
rect 11431 -3897 11487 -3888
rect 11431 -3962 11487 -3953
rect 12599 -3897 12655 -3888
rect 12599 -3962 12655 -3953
rect 13767 -3897 13823 -3888
rect 13767 -3962 13823 -3953
rect 14935 -3897 14991 -3888
rect 14935 -3962 14991 -3953
rect 16103 -3897 16159 -3888
rect 16103 -3962 16159 -3953
rect 17271 -3897 17327 -3888
rect 17271 -3962 17327 -3953
rect 18439 -3897 18495 -3888
rect 18439 -3962 18495 -3953
rect 19607 -3897 19663 -3888
rect 19607 -3962 19663 -3953
rect 20775 -3897 20831 -3888
rect 20775 -3962 20831 -3953
rect 21943 -3897 21999 -3888
rect 21943 -3962 21999 -3953
rect 23111 -3897 23167 -3888
rect 23111 -3962 23167 -3953
rect 24279 -3897 24335 -3888
rect 24279 -3962 24335 -3953
rect 25447 -3897 25503 -3888
rect 25447 -3962 25503 -3953
rect 26615 -3897 26671 -3888
rect 26615 -3962 26671 -3953
rect 27783 -3897 27839 -3888
rect 27783 -3962 27839 -3953
rect 28951 -3897 29007 -3888
rect 28951 -3962 29007 -3953
rect 30119 -3897 30175 -3888
rect 30119 -3962 30175 -3953
rect 31287 -3897 31343 -3888
rect 31287 -3962 31343 -3953
rect 32455 -3897 32511 -3888
rect 32455 -3962 32511 -3953
rect 33623 -3897 33679 -3888
rect 33623 -3962 33679 -3953
rect 34791 -3897 34847 -3888
rect 34791 -3962 34847 -3953
rect 35959 -3897 36015 -3888
rect 35959 -3962 36015 -3953
rect 37127 -3897 37183 -3888
rect 37127 -3962 37183 -3953
rect 38295 -3897 38351 -3888
rect 38295 -3962 38351 -3953
rect 39463 -3897 39519 -3888
rect 39463 -3962 39519 -3953
rect 40631 -3897 40687 -3888
rect 40631 -3962 40687 -3953
rect 41799 -3897 41855 -3888
rect 41799 -3962 41855 -3953
rect 42967 -3897 43023 -3888
rect 42967 -3962 43023 -3953
rect 44135 -3897 44191 -3888
rect 44135 -3962 44191 -3953
<< via2 >>
rect 13914 1451 13970 1453
rect 13914 1399 13916 1451
rect 13916 1399 13968 1451
rect 13968 1399 13970 1451
rect 13914 1397 13970 1399
rect 15162 1451 15218 1453
rect 15162 1399 15164 1451
rect 15164 1399 15216 1451
rect 15216 1399 15218 1451
rect 15162 1397 15218 1399
rect 16410 1451 16466 1453
rect 16410 1399 16412 1451
rect 16412 1399 16464 1451
rect 16464 1399 16466 1451
rect 16410 1397 16466 1399
rect 17658 1451 17714 1453
rect 17658 1399 17660 1451
rect 17660 1399 17712 1451
rect 17712 1399 17714 1451
rect 17658 1397 17714 1399
rect 18906 1451 18962 1453
rect 18906 1399 18908 1451
rect 18908 1399 18960 1451
rect 18960 1399 18962 1451
rect 18906 1397 18962 1399
rect 20154 1451 20210 1453
rect 20154 1399 20156 1451
rect 20156 1399 20208 1451
rect 20208 1399 20210 1451
rect 20154 1397 20210 1399
rect 21402 1451 21458 1453
rect 21402 1399 21404 1451
rect 21404 1399 21456 1451
rect 21456 1399 21458 1451
rect 21402 1397 21458 1399
rect 22650 1451 22706 1453
rect 22650 1399 22652 1451
rect 22652 1399 22704 1451
rect 22704 1399 22706 1451
rect 22650 1397 22706 1399
rect 23898 1451 23954 1453
rect 23898 1399 23900 1451
rect 23900 1399 23952 1451
rect 23952 1399 23954 1451
rect 23898 1397 23954 1399
rect 25146 1451 25202 1453
rect 25146 1399 25148 1451
rect 25148 1399 25200 1451
rect 25200 1399 25202 1451
rect 25146 1397 25202 1399
rect 26394 1451 26450 1453
rect 26394 1399 26396 1451
rect 26396 1399 26448 1451
rect 26448 1399 26450 1451
rect 26394 1397 26450 1399
rect 27642 1451 27698 1453
rect 27642 1399 27644 1451
rect 27644 1399 27696 1451
rect 27696 1399 27698 1451
rect 27642 1397 27698 1399
rect 28890 1451 28946 1453
rect 28890 1399 28892 1451
rect 28892 1399 28944 1451
rect 28944 1399 28946 1451
rect 28890 1397 28946 1399
rect 30138 1451 30194 1453
rect 30138 1399 30140 1451
rect 30140 1399 30192 1451
rect 30192 1399 30194 1451
rect 30138 1397 30194 1399
rect 31386 1451 31442 1453
rect 31386 1399 31388 1451
rect 31388 1399 31440 1451
rect 31440 1399 31442 1451
rect 31386 1397 31442 1399
rect 32634 1451 32690 1453
rect 32634 1399 32636 1451
rect 32636 1399 32688 1451
rect 32688 1399 32690 1451
rect 32634 1397 32690 1399
rect 33882 1451 33938 1453
rect 33882 1399 33884 1451
rect 33884 1399 33936 1451
rect 33936 1399 33938 1451
rect 33882 1397 33938 1399
rect 35130 1451 35186 1453
rect 35130 1399 35132 1451
rect 35132 1399 35184 1451
rect 35184 1399 35186 1451
rect 35130 1397 35186 1399
rect 36378 1451 36434 1453
rect 36378 1399 36380 1451
rect 36380 1399 36432 1451
rect 36432 1399 36434 1451
rect 36378 1397 36434 1399
rect 37626 1451 37682 1453
rect 37626 1399 37628 1451
rect 37628 1399 37680 1451
rect 37680 1399 37682 1451
rect 37626 1397 37682 1399
rect 38874 1451 38930 1453
rect 38874 1399 38876 1451
rect 38876 1399 38928 1451
rect 38928 1399 38930 1451
rect 38874 1397 38930 1399
rect 40122 1451 40178 1453
rect 40122 1399 40124 1451
rect 40124 1399 40176 1451
rect 40176 1399 40178 1451
rect 40122 1397 40178 1399
rect 41370 1451 41426 1453
rect 41370 1399 41372 1451
rect 41372 1399 41424 1451
rect 41424 1399 41426 1451
rect 41370 1397 41426 1399
rect 42618 1451 42674 1453
rect 42618 1399 42620 1451
rect 42620 1399 42672 1451
rect 42672 1399 42674 1451
rect 42618 1397 42674 1399
rect 43866 1451 43922 1453
rect 43866 1399 43868 1451
rect 43868 1399 43920 1451
rect 43920 1399 43922 1451
rect 43866 1397 43922 1399
rect 45114 1451 45170 1453
rect 45114 1399 45116 1451
rect 45116 1399 45168 1451
rect 45168 1399 45170 1451
rect 45114 1397 45170 1399
rect 46362 1451 46418 1453
rect 46362 1399 46364 1451
rect 46364 1399 46416 1451
rect 46416 1399 46418 1451
rect 46362 1397 46418 1399
rect 47610 1451 47666 1453
rect 47610 1399 47612 1451
rect 47612 1399 47664 1451
rect 47664 1399 47666 1451
rect 47610 1397 47666 1399
rect 48858 1451 48914 1453
rect 48858 1399 48860 1451
rect 48860 1399 48912 1451
rect 48912 1399 48914 1451
rect 48858 1397 48914 1399
rect 50106 1451 50162 1453
rect 50106 1399 50108 1451
rect 50108 1399 50160 1451
rect 50160 1399 50162 1451
rect 50106 1397 50162 1399
rect 51354 1451 51410 1453
rect 51354 1399 51356 1451
rect 51356 1399 51408 1451
rect 51408 1399 51410 1451
rect 51354 1397 51410 1399
rect 52602 1451 52658 1453
rect 52602 1399 52604 1451
rect 52604 1399 52656 1451
rect 52656 1399 52658 1451
rect 52602 1397 52658 1399
rect 13629 277 13685 333
rect 23613 277 23669 333
rect 33597 277 33653 333
rect 43581 277 43637 333
rect 3255 -3953 3311 -3897
rect 4423 -3953 4479 -3897
rect 5591 -3953 5647 -3897
rect 6759 -3953 6815 -3897
rect 7927 -3953 7983 -3897
rect 9095 -3953 9151 -3897
rect 10263 -3953 10319 -3897
rect 11431 -3953 11487 -3897
rect 12599 -3953 12655 -3897
rect 13767 -3953 13823 -3897
rect 14935 -3953 14991 -3897
rect 16103 -3953 16159 -3897
rect 17271 -3953 17327 -3897
rect 18439 -3953 18495 -3897
rect 19607 -3953 19663 -3897
rect 20775 -3953 20831 -3897
rect 21943 -3953 21999 -3897
rect 23111 -3953 23167 -3897
rect 24279 -3953 24335 -3897
rect 25447 -3953 25503 -3897
rect 26615 -3953 26671 -3897
rect 27783 -3953 27839 -3897
rect 28951 -3953 29007 -3897
rect 30119 -3953 30175 -3897
rect 31287 -3953 31343 -3897
rect 32455 -3953 32511 -3897
rect 33623 -3953 33679 -3897
rect 34791 -3953 34847 -3897
rect 35959 -3953 36015 -3897
rect 37127 -3953 37183 -3897
rect 38295 -3953 38351 -3897
rect 39463 -3953 39519 -3897
rect 40631 -3953 40687 -3897
rect 41799 -3953 41855 -3897
rect 42967 -3953 43023 -3897
rect 44135 -3953 44191 -3897
<< metal3 >>
rect 13909 1457 13975 1458
rect 15157 1457 15223 1458
rect 16405 1457 16471 1458
rect 17653 1457 17719 1458
rect 18901 1457 18967 1458
rect 20149 1457 20215 1458
rect 21397 1457 21463 1458
rect 22645 1457 22711 1458
rect 23893 1457 23959 1458
rect 25141 1457 25207 1458
rect 26389 1457 26455 1458
rect 27637 1457 27703 1458
rect 28885 1457 28951 1458
rect 30133 1457 30199 1458
rect 31381 1457 31447 1458
rect 32629 1457 32695 1458
rect 33877 1457 33943 1458
rect 35125 1457 35191 1458
rect 36373 1457 36439 1458
rect 37621 1457 37687 1458
rect 38869 1457 38935 1458
rect 40117 1457 40183 1458
rect 41365 1457 41431 1458
rect 42613 1457 42679 1458
rect 43861 1457 43927 1458
rect 45109 1457 45175 1458
rect 46357 1457 46423 1458
rect 47605 1457 47671 1458
rect 48853 1457 48919 1458
rect 50101 1457 50167 1458
rect 51349 1457 51415 1458
rect 52597 1457 52663 1458
rect 13867 1393 13910 1457
rect 13974 1393 14017 1457
rect 15115 1393 15158 1457
rect 15222 1393 15265 1457
rect 16363 1393 16406 1457
rect 16470 1393 16513 1457
rect 17611 1393 17654 1457
rect 17718 1393 17761 1457
rect 18859 1393 18902 1457
rect 18966 1393 19009 1457
rect 20107 1393 20150 1457
rect 20214 1393 20257 1457
rect 21355 1393 21398 1457
rect 21462 1393 21505 1457
rect 22603 1393 22646 1457
rect 22710 1393 22753 1457
rect 23851 1393 23894 1457
rect 23958 1393 24001 1457
rect 25099 1393 25142 1457
rect 25206 1393 25249 1457
rect 26347 1393 26390 1457
rect 26454 1393 26497 1457
rect 27595 1393 27638 1457
rect 27702 1393 27745 1457
rect 28843 1393 28886 1457
rect 28950 1393 28993 1457
rect 30091 1393 30134 1457
rect 30198 1393 30241 1457
rect 31339 1393 31382 1457
rect 31446 1393 31489 1457
rect 32587 1393 32630 1457
rect 32694 1393 32737 1457
rect 33835 1393 33878 1457
rect 33942 1393 33985 1457
rect 35083 1393 35126 1457
rect 35190 1393 35233 1457
rect 36331 1393 36374 1457
rect 36438 1393 36481 1457
rect 37579 1393 37622 1457
rect 37686 1393 37729 1457
rect 38827 1393 38870 1457
rect 38934 1393 38977 1457
rect 40075 1393 40118 1457
rect 40182 1393 40225 1457
rect 41323 1393 41366 1457
rect 41430 1393 41473 1457
rect 42571 1393 42614 1457
rect 42678 1393 42721 1457
rect 43819 1393 43862 1457
rect 43926 1393 43969 1457
rect 45067 1393 45110 1457
rect 45174 1393 45217 1457
rect 46315 1393 46358 1457
rect 46422 1393 46465 1457
rect 47563 1393 47606 1457
rect 47670 1393 47713 1457
rect 48811 1393 48854 1457
rect 48918 1393 48961 1457
rect 50059 1393 50102 1457
rect 50166 1393 50209 1457
rect 51307 1393 51350 1457
rect 51414 1393 51457 1457
rect 52555 1393 52598 1457
rect 52662 1393 52705 1457
rect 13909 1392 13975 1393
rect 15157 1392 15223 1393
rect 16405 1392 16471 1393
rect 17653 1392 17719 1393
rect 18901 1392 18967 1393
rect 20149 1392 20215 1393
rect 21397 1392 21463 1393
rect 22645 1392 22711 1393
rect 23893 1392 23959 1393
rect 25141 1392 25207 1393
rect 26389 1392 26455 1393
rect 27637 1392 27703 1393
rect 28885 1392 28951 1393
rect 30133 1392 30199 1393
rect 31381 1392 31447 1393
rect 32629 1392 32695 1393
rect 33877 1392 33943 1393
rect 35125 1392 35191 1393
rect 36373 1392 36439 1393
rect 37621 1392 37687 1393
rect 38869 1392 38935 1393
rect 40117 1392 40183 1393
rect 41365 1392 41431 1393
rect 42613 1392 42679 1393
rect 43861 1392 43927 1393
rect 45109 1392 45175 1393
rect 46357 1392 46423 1393
rect 47605 1392 47671 1393
rect 48853 1392 48919 1393
rect 50101 1392 50167 1393
rect 51349 1392 51415 1393
rect 52597 1392 52663 1393
rect 13624 337 13690 338
rect 23608 337 23674 338
rect 33592 337 33658 338
rect 43576 337 43642 338
rect 13582 273 13625 337
rect 13689 273 13732 337
rect 23566 273 23609 337
rect 23673 273 23716 337
rect 33550 273 33593 337
rect 33657 273 33700 337
rect 43534 273 43577 337
rect 43641 273 43684 337
rect 13624 272 13690 273
rect 23608 272 23674 273
rect 33592 272 33658 273
rect 43576 272 43642 273
rect 25437 -516 25443 -452
rect 25507 -454 25513 -452
rect 32624 -454 32630 -452
rect 25507 -514 32630 -454
rect 25507 -516 25513 -514
rect 32624 -516 32630 -514
rect 32694 -516 32700 -452
rect 9085 -760 9091 -696
rect 9155 -698 9161 -696
rect 15152 -698 15158 -696
rect 9155 -758 15158 -698
rect 9155 -760 9161 -758
rect 15152 -760 15158 -758
rect 15222 -760 15228 -696
rect 24269 -760 24275 -696
rect 24339 -698 24345 -696
rect 31376 -698 31382 -696
rect 24339 -758 31382 -698
rect 24339 -760 24345 -758
rect 31376 -760 31382 -758
rect 31446 -760 31452 -696
rect 5581 -1004 5587 -940
rect 5651 -942 5657 -940
rect 33587 -942 33593 -940
rect 5651 -1002 33593 -942
rect 5651 -1004 5657 -1002
rect 33587 -1004 33593 -1002
rect 33657 -1004 33663 -940
rect 7917 -1248 7923 -1184
rect 7987 -1186 7993 -1184
rect 13904 -1186 13910 -1184
rect 7987 -1246 13910 -1186
rect 7987 -1248 7993 -1246
rect 13904 -1248 13910 -1246
rect 13974 -1248 13980 -1184
rect 16093 -1248 16099 -1184
rect 16163 -1186 16169 -1184
rect 22640 -1186 22646 -1184
rect 16163 -1246 22646 -1186
rect 16163 -1248 16169 -1246
rect 22640 -1248 22646 -1246
rect 22710 -1248 22716 -1184
rect 23101 -1248 23107 -1184
rect 23171 -1186 23177 -1184
rect 30128 -1186 30134 -1184
rect 23171 -1246 30134 -1186
rect 23171 -1248 23177 -1246
rect 30128 -1248 30134 -1246
rect 30198 -1248 30204 -1184
rect 33613 -1248 33619 -1184
rect 33683 -1186 33689 -1184
rect 41360 -1186 41366 -1184
rect 33683 -1246 41366 -1186
rect 33683 -1248 33689 -1246
rect 41360 -1248 41366 -1246
rect 41430 -1248 41436 -1184
rect 41789 -1248 41795 -1184
rect 41859 -1186 41865 -1184
rect 50096 -1186 50102 -1184
rect 41859 -1246 50102 -1186
rect 41859 -1248 41865 -1246
rect 50096 -1248 50102 -1246
rect 50166 -1248 50172 -1184
rect 3245 -1492 3251 -1428
rect 3315 -1430 3321 -1428
rect 13619 -1430 13625 -1428
rect 3315 -1490 13625 -1430
rect 3315 -1492 3321 -1490
rect 13619 -1492 13625 -1490
rect 13689 -1492 13695 -1428
rect 14925 -1492 14931 -1428
rect 14995 -1430 15001 -1428
rect 21392 -1430 21398 -1428
rect 14995 -1490 21398 -1430
rect 14995 -1492 15001 -1490
rect 21392 -1492 21398 -1490
rect 21462 -1492 21468 -1428
rect 21933 -1492 21939 -1428
rect 22003 -1430 22009 -1428
rect 28880 -1430 28886 -1428
rect 22003 -1490 28886 -1430
rect 22003 -1492 22009 -1490
rect 28880 -1492 28886 -1490
rect 28950 -1492 28956 -1428
rect 32445 -1492 32451 -1428
rect 32515 -1430 32521 -1428
rect 40112 -1430 40118 -1428
rect 32515 -1490 40118 -1430
rect 32515 -1492 32521 -1490
rect 40112 -1492 40118 -1490
rect 40182 -1492 40188 -1428
rect 40621 -1492 40627 -1428
rect 40691 -1430 40697 -1428
rect 48848 -1430 48854 -1428
rect 40691 -1490 48854 -1430
rect 40691 -1492 40697 -1490
rect 48848 -1492 48854 -1490
rect 48918 -1492 48924 -1428
rect 13757 -1736 13763 -1672
rect 13827 -1674 13833 -1672
rect 20144 -1674 20150 -1672
rect 13827 -1734 20150 -1674
rect 13827 -1736 13833 -1734
rect 20144 -1736 20150 -1734
rect 20214 -1736 20220 -1672
rect 20765 -1736 20771 -1672
rect 20835 -1674 20841 -1672
rect 27632 -1674 27638 -1672
rect 20835 -1734 27638 -1674
rect 20835 -1736 20841 -1734
rect 27632 -1736 27638 -1734
rect 27702 -1736 27708 -1672
rect 31277 -1736 31283 -1672
rect 31347 -1674 31353 -1672
rect 38864 -1674 38870 -1672
rect 31347 -1734 38870 -1674
rect 31347 -1736 31353 -1734
rect 38864 -1736 38870 -1734
rect 38934 -1736 38940 -1672
rect 39453 -1736 39459 -1672
rect 39523 -1674 39529 -1672
rect 47600 -1674 47606 -1672
rect 39523 -1734 47606 -1674
rect 39523 -1736 39529 -1734
rect 47600 -1736 47606 -1734
rect 47670 -1736 47676 -1672
rect 12589 -1980 12595 -1916
rect 12659 -1918 12665 -1916
rect 18896 -1918 18902 -1916
rect 12659 -1978 18902 -1918
rect 12659 -1980 12665 -1978
rect 18896 -1980 18902 -1978
rect 18966 -1980 18972 -1916
rect 19597 -1980 19603 -1916
rect 19667 -1918 19673 -1916
rect 26384 -1918 26390 -1916
rect 19667 -1978 26390 -1918
rect 19667 -1980 19673 -1978
rect 26384 -1980 26390 -1978
rect 26454 -1980 26460 -1916
rect 30109 -1980 30115 -1916
rect 30179 -1918 30185 -1916
rect 37616 -1918 37622 -1916
rect 30179 -1978 37622 -1918
rect 30179 -1980 30185 -1978
rect 37616 -1980 37622 -1978
rect 37686 -1980 37692 -1916
rect 38285 -1980 38291 -1916
rect 38355 -1918 38361 -1916
rect 46352 -1918 46358 -1916
rect 38355 -1978 46358 -1918
rect 38355 -1980 38361 -1978
rect 46352 -1980 46358 -1978
rect 46422 -1980 46428 -1916
rect 11421 -2224 11427 -2160
rect 11491 -2162 11497 -2160
rect 17648 -2162 17654 -2160
rect 11491 -2222 17654 -2162
rect 11491 -2224 11497 -2222
rect 17648 -2224 17654 -2222
rect 17718 -2224 17724 -2160
rect 18429 -2224 18435 -2160
rect 18499 -2162 18505 -2160
rect 25136 -2162 25142 -2160
rect 18499 -2222 25142 -2162
rect 18499 -2224 18505 -2222
rect 25136 -2224 25142 -2222
rect 25206 -2224 25212 -2160
rect 28941 -2224 28947 -2160
rect 29011 -2162 29017 -2160
rect 36368 -2162 36374 -2160
rect 29011 -2222 36374 -2162
rect 29011 -2224 29017 -2222
rect 36368 -2224 36374 -2222
rect 36438 -2224 36444 -2160
rect 37117 -2224 37123 -2160
rect 37187 -2162 37193 -2160
rect 45104 -2162 45110 -2160
rect 37187 -2222 45110 -2162
rect 37187 -2224 37193 -2222
rect 45104 -2224 45110 -2222
rect 45174 -2224 45180 -2160
rect 10253 -2468 10259 -2404
rect 10323 -2406 10329 -2404
rect 16400 -2406 16406 -2404
rect 10323 -2466 16406 -2406
rect 10323 -2468 10329 -2466
rect 16400 -2468 16406 -2466
rect 16470 -2468 16476 -2404
rect 17261 -2468 17267 -2404
rect 17331 -2406 17337 -2404
rect 23888 -2406 23894 -2404
rect 17331 -2466 23894 -2406
rect 17331 -2468 17337 -2466
rect 23888 -2468 23894 -2466
rect 23958 -2468 23964 -2404
rect 27773 -2468 27779 -2404
rect 27843 -2406 27849 -2404
rect 35120 -2406 35126 -2404
rect 27843 -2466 35126 -2406
rect 27843 -2468 27849 -2466
rect 35120 -2468 35126 -2466
rect 35190 -2468 35196 -2404
rect 35949 -2468 35955 -2404
rect 36019 -2406 36025 -2404
rect 43856 -2406 43862 -2404
rect 36019 -2466 43862 -2406
rect 36019 -2468 36025 -2466
rect 43856 -2468 43862 -2466
rect 43926 -2468 43932 -2404
rect 6749 -2712 6755 -2648
rect 6819 -2650 6825 -2648
rect 43571 -2650 43577 -2648
rect 6819 -2710 43577 -2650
rect 6819 -2712 6825 -2710
rect 43571 -2712 43577 -2710
rect 43641 -2712 43647 -2648
rect 44125 -2712 44131 -2648
rect 44195 -2650 44201 -2648
rect 52592 -2650 52598 -2648
rect 44195 -2710 52598 -2650
rect 44195 -2712 44201 -2710
rect 52592 -2712 52598 -2710
rect 52662 -2712 52668 -2648
rect 4413 -2956 4419 -2892
rect 4483 -2894 4489 -2892
rect 23603 -2894 23609 -2892
rect 4483 -2954 23609 -2894
rect 4483 -2956 4489 -2954
rect 23603 -2956 23609 -2954
rect 23673 -2956 23679 -2892
rect 26605 -2956 26611 -2892
rect 26675 -2894 26681 -2892
rect 33872 -2894 33878 -2892
rect 26675 -2954 33878 -2894
rect 26675 -2956 26681 -2954
rect 33872 -2956 33878 -2954
rect 33942 -2956 33948 -2892
rect 34781 -2956 34787 -2892
rect 34851 -2894 34857 -2892
rect 42608 -2894 42614 -2892
rect 34851 -2954 42614 -2894
rect 34851 -2956 34857 -2954
rect 42608 -2956 42614 -2954
rect 42678 -2956 42684 -2892
rect 42957 -2956 42963 -2892
rect 43027 -2894 43033 -2892
rect 51344 -2894 51350 -2892
rect 43027 -2954 51350 -2894
rect 43027 -2956 43033 -2954
rect 51344 -2956 51350 -2954
rect 51414 -2956 51420 -2892
rect 3250 -3893 3316 -3892
rect 4418 -3893 4484 -3892
rect 5586 -3893 5652 -3892
rect 6754 -3893 6820 -3892
rect 7922 -3893 7988 -3892
rect 9090 -3893 9156 -3892
rect 10258 -3893 10324 -3892
rect 11426 -3893 11492 -3892
rect 12594 -3893 12660 -3892
rect 13762 -3893 13828 -3892
rect 14930 -3893 14996 -3892
rect 16098 -3893 16164 -3892
rect 17266 -3893 17332 -3892
rect 18434 -3893 18500 -3892
rect 19602 -3893 19668 -3892
rect 20770 -3893 20836 -3892
rect 21938 -3893 22004 -3892
rect 23106 -3893 23172 -3892
rect 24274 -3893 24340 -3892
rect 25442 -3893 25508 -3892
rect 26610 -3893 26676 -3892
rect 27778 -3893 27844 -3892
rect 28946 -3893 29012 -3892
rect 30114 -3893 30180 -3892
rect 31282 -3893 31348 -3892
rect 32450 -3893 32516 -3892
rect 33618 -3893 33684 -3892
rect 34786 -3893 34852 -3892
rect 35954 -3893 36020 -3892
rect 37122 -3893 37188 -3892
rect 38290 -3893 38356 -3892
rect 39458 -3893 39524 -3892
rect 40626 -3893 40692 -3892
rect 41794 -3893 41860 -3892
rect 42962 -3893 43028 -3892
rect 44130 -3893 44196 -3892
rect 3208 -3957 3251 -3893
rect 3315 -3957 3358 -3893
rect 4376 -3957 4419 -3893
rect 4483 -3957 4526 -3893
rect 5544 -3957 5587 -3893
rect 5651 -3957 5694 -3893
rect 6712 -3957 6755 -3893
rect 6819 -3957 6862 -3893
rect 7880 -3957 7923 -3893
rect 7987 -3957 8030 -3893
rect 9048 -3957 9091 -3893
rect 9155 -3957 9198 -3893
rect 10216 -3957 10259 -3893
rect 10323 -3957 10366 -3893
rect 11384 -3957 11427 -3893
rect 11491 -3957 11534 -3893
rect 12552 -3957 12595 -3893
rect 12659 -3957 12702 -3893
rect 13720 -3957 13763 -3893
rect 13827 -3957 13870 -3893
rect 14888 -3957 14931 -3893
rect 14995 -3957 15038 -3893
rect 16056 -3957 16099 -3893
rect 16163 -3957 16206 -3893
rect 17224 -3957 17267 -3893
rect 17331 -3957 17374 -3893
rect 18392 -3957 18435 -3893
rect 18499 -3957 18542 -3893
rect 19560 -3957 19603 -3893
rect 19667 -3957 19710 -3893
rect 20728 -3957 20771 -3893
rect 20835 -3957 20878 -3893
rect 21896 -3957 21939 -3893
rect 22003 -3957 22046 -3893
rect 23064 -3957 23107 -3893
rect 23171 -3957 23214 -3893
rect 24232 -3957 24275 -3893
rect 24339 -3957 24382 -3893
rect 25400 -3957 25443 -3893
rect 25507 -3957 25550 -3893
rect 26568 -3957 26611 -3893
rect 26675 -3957 26718 -3893
rect 27736 -3957 27779 -3893
rect 27843 -3957 27886 -3893
rect 28904 -3957 28947 -3893
rect 29011 -3957 29054 -3893
rect 30072 -3957 30115 -3893
rect 30179 -3957 30222 -3893
rect 31240 -3957 31283 -3893
rect 31347 -3957 31390 -3893
rect 32408 -3957 32451 -3893
rect 32515 -3957 32558 -3893
rect 33576 -3957 33619 -3893
rect 33683 -3957 33726 -3893
rect 34744 -3957 34787 -3893
rect 34851 -3957 34894 -3893
rect 35912 -3957 35955 -3893
rect 36019 -3957 36062 -3893
rect 37080 -3957 37123 -3893
rect 37187 -3957 37230 -3893
rect 38248 -3957 38291 -3893
rect 38355 -3957 38398 -3893
rect 39416 -3957 39459 -3893
rect 39523 -3957 39566 -3893
rect 40584 -3957 40627 -3893
rect 40691 -3957 40734 -3893
rect 41752 -3957 41795 -3893
rect 41859 -3957 41902 -3893
rect 42920 -3957 42963 -3893
rect 43027 -3957 43070 -3893
rect 44088 -3957 44131 -3893
rect 44195 -3957 44238 -3893
rect 3250 -3958 3316 -3957
rect 4418 -3958 4484 -3957
rect 5586 -3958 5652 -3957
rect 6754 -3958 6820 -3957
rect 7922 -3958 7988 -3957
rect 9090 -3958 9156 -3957
rect 10258 -3958 10324 -3957
rect 11426 -3958 11492 -3957
rect 12594 -3958 12660 -3957
rect 13762 -3958 13828 -3957
rect 14930 -3958 14996 -3957
rect 16098 -3958 16164 -3957
rect 17266 -3958 17332 -3957
rect 18434 -3958 18500 -3957
rect 19602 -3958 19668 -3957
rect 20770 -3958 20836 -3957
rect 21938 -3958 22004 -3957
rect 23106 -3958 23172 -3957
rect 24274 -3958 24340 -3957
rect 25442 -3958 25508 -3957
rect 26610 -3958 26676 -3957
rect 27778 -3958 27844 -3957
rect 28946 -3958 29012 -3957
rect 30114 -3958 30180 -3957
rect 31282 -3958 31348 -3957
rect 32450 -3958 32516 -3957
rect 33618 -3958 33684 -3957
rect 34786 -3958 34852 -3957
rect 35954 -3958 36020 -3957
rect 37122 -3958 37188 -3957
rect 38290 -3958 38356 -3957
rect 39458 -3958 39524 -3957
rect 40626 -3958 40692 -3957
rect 41794 -3958 41860 -3957
rect 42962 -3958 43028 -3957
rect 44130 -3958 44196 -3957
<< via3 >>
rect 13910 1453 13974 1457
rect 13910 1397 13914 1453
rect 13914 1397 13970 1453
rect 13970 1397 13974 1453
rect 13910 1393 13974 1397
rect 15158 1453 15222 1457
rect 15158 1397 15162 1453
rect 15162 1397 15218 1453
rect 15218 1397 15222 1453
rect 15158 1393 15222 1397
rect 16406 1453 16470 1457
rect 16406 1397 16410 1453
rect 16410 1397 16466 1453
rect 16466 1397 16470 1453
rect 16406 1393 16470 1397
rect 17654 1453 17718 1457
rect 17654 1397 17658 1453
rect 17658 1397 17714 1453
rect 17714 1397 17718 1453
rect 17654 1393 17718 1397
rect 18902 1453 18966 1457
rect 18902 1397 18906 1453
rect 18906 1397 18962 1453
rect 18962 1397 18966 1453
rect 18902 1393 18966 1397
rect 20150 1453 20214 1457
rect 20150 1397 20154 1453
rect 20154 1397 20210 1453
rect 20210 1397 20214 1453
rect 20150 1393 20214 1397
rect 21398 1453 21462 1457
rect 21398 1397 21402 1453
rect 21402 1397 21458 1453
rect 21458 1397 21462 1453
rect 21398 1393 21462 1397
rect 22646 1453 22710 1457
rect 22646 1397 22650 1453
rect 22650 1397 22706 1453
rect 22706 1397 22710 1453
rect 22646 1393 22710 1397
rect 23894 1453 23958 1457
rect 23894 1397 23898 1453
rect 23898 1397 23954 1453
rect 23954 1397 23958 1453
rect 23894 1393 23958 1397
rect 25142 1453 25206 1457
rect 25142 1397 25146 1453
rect 25146 1397 25202 1453
rect 25202 1397 25206 1453
rect 25142 1393 25206 1397
rect 26390 1453 26454 1457
rect 26390 1397 26394 1453
rect 26394 1397 26450 1453
rect 26450 1397 26454 1453
rect 26390 1393 26454 1397
rect 27638 1453 27702 1457
rect 27638 1397 27642 1453
rect 27642 1397 27698 1453
rect 27698 1397 27702 1453
rect 27638 1393 27702 1397
rect 28886 1453 28950 1457
rect 28886 1397 28890 1453
rect 28890 1397 28946 1453
rect 28946 1397 28950 1453
rect 28886 1393 28950 1397
rect 30134 1453 30198 1457
rect 30134 1397 30138 1453
rect 30138 1397 30194 1453
rect 30194 1397 30198 1453
rect 30134 1393 30198 1397
rect 31382 1453 31446 1457
rect 31382 1397 31386 1453
rect 31386 1397 31442 1453
rect 31442 1397 31446 1453
rect 31382 1393 31446 1397
rect 32630 1453 32694 1457
rect 32630 1397 32634 1453
rect 32634 1397 32690 1453
rect 32690 1397 32694 1453
rect 32630 1393 32694 1397
rect 33878 1453 33942 1457
rect 33878 1397 33882 1453
rect 33882 1397 33938 1453
rect 33938 1397 33942 1453
rect 33878 1393 33942 1397
rect 35126 1453 35190 1457
rect 35126 1397 35130 1453
rect 35130 1397 35186 1453
rect 35186 1397 35190 1453
rect 35126 1393 35190 1397
rect 36374 1453 36438 1457
rect 36374 1397 36378 1453
rect 36378 1397 36434 1453
rect 36434 1397 36438 1453
rect 36374 1393 36438 1397
rect 37622 1453 37686 1457
rect 37622 1397 37626 1453
rect 37626 1397 37682 1453
rect 37682 1397 37686 1453
rect 37622 1393 37686 1397
rect 38870 1453 38934 1457
rect 38870 1397 38874 1453
rect 38874 1397 38930 1453
rect 38930 1397 38934 1453
rect 38870 1393 38934 1397
rect 40118 1453 40182 1457
rect 40118 1397 40122 1453
rect 40122 1397 40178 1453
rect 40178 1397 40182 1453
rect 40118 1393 40182 1397
rect 41366 1453 41430 1457
rect 41366 1397 41370 1453
rect 41370 1397 41426 1453
rect 41426 1397 41430 1453
rect 41366 1393 41430 1397
rect 42614 1453 42678 1457
rect 42614 1397 42618 1453
rect 42618 1397 42674 1453
rect 42674 1397 42678 1453
rect 42614 1393 42678 1397
rect 43862 1453 43926 1457
rect 43862 1397 43866 1453
rect 43866 1397 43922 1453
rect 43922 1397 43926 1453
rect 43862 1393 43926 1397
rect 45110 1453 45174 1457
rect 45110 1397 45114 1453
rect 45114 1397 45170 1453
rect 45170 1397 45174 1453
rect 45110 1393 45174 1397
rect 46358 1453 46422 1457
rect 46358 1397 46362 1453
rect 46362 1397 46418 1453
rect 46418 1397 46422 1453
rect 46358 1393 46422 1397
rect 47606 1453 47670 1457
rect 47606 1397 47610 1453
rect 47610 1397 47666 1453
rect 47666 1397 47670 1453
rect 47606 1393 47670 1397
rect 48854 1453 48918 1457
rect 48854 1397 48858 1453
rect 48858 1397 48914 1453
rect 48914 1397 48918 1453
rect 48854 1393 48918 1397
rect 50102 1453 50166 1457
rect 50102 1397 50106 1453
rect 50106 1397 50162 1453
rect 50162 1397 50166 1453
rect 50102 1393 50166 1397
rect 51350 1453 51414 1457
rect 51350 1397 51354 1453
rect 51354 1397 51410 1453
rect 51410 1397 51414 1453
rect 51350 1393 51414 1397
rect 52598 1453 52662 1457
rect 52598 1397 52602 1453
rect 52602 1397 52658 1453
rect 52658 1397 52662 1453
rect 52598 1393 52662 1397
rect 13625 333 13689 337
rect 13625 277 13629 333
rect 13629 277 13685 333
rect 13685 277 13689 333
rect 13625 273 13689 277
rect 23609 333 23673 337
rect 23609 277 23613 333
rect 23613 277 23669 333
rect 23669 277 23673 333
rect 23609 273 23673 277
rect 33593 333 33657 337
rect 33593 277 33597 333
rect 33597 277 33653 333
rect 33653 277 33657 333
rect 33593 273 33657 277
rect 43577 333 43641 337
rect 43577 277 43581 333
rect 43581 277 43637 333
rect 43637 277 43641 333
rect 43577 273 43641 277
rect 25443 -516 25507 -452
rect 32630 -516 32694 -452
rect 9091 -760 9155 -696
rect 15158 -760 15222 -696
rect 24275 -760 24339 -696
rect 31382 -760 31446 -696
rect 5587 -1004 5651 -940
rect 33593 -1004 33657 -940
rect 7923 -1248 7987 -1184
rect 13910 -1248 13974 -1184
rect 16099 -1248 16163 -1184
rect 22646 -1248 22710 -1184
rect 23107 -1248 23171 -1184
rect 30134 -1248 30198 -1184
rect 33619 -1248 33683 -1184
rect 41366 -1248 41430 -1184
rect 41795 -1248 41859 -1184
rect 50102 -1248 50166 -1184
rect 3251 -1492 3315 -1428
rect 13625 -1492 13689 -1428
rect 14931 -1492 14995 -1428
rect 21398 -1492 21462 -1428
rect 21939 -1492 22003 -1428
rect 28886 -1492 28950 -1428
rect 32451 -1492 32515 -1428
rect 40118 -1492 40182 -1428
rect 40627 -1492 40691 -1428
rect 48854 -1492 48918 -1428
rect 13763 -1736 13827 -1672
rect 20150 -1736 20214 -1672
rect 20771 -1736 20835 -1672
rect 27638 -1736 27702 -1672
rect 31283 -1736 31347 -1672
rect 38870 -1736 38934 -1672
rect 39459 -1736 39523 -1672
rect 47606 -1736 47670 -1672
rect 12595 -1980 12659 -1916
rect 18902 -1980 18966 -1916
rect 19603 -1980 19667 -1916
rect 26390 -1980 26454 -1916
rect 30115 -1980 30179 -1916
rect 37622 -1980 37686 -1916
rect 38291 -1980 38355 -1916
rect 46358 -1980 46422 -1916
rect 11427 -2224 11491 -2160
rect 17654 -2224 17718 -2160
rect 18435 -2224 18499 -2160
rect 25142 -2224 25206 -2160
rect 28947 -2224 29011 -2160
rect 36374 -2224 36438 -2160
rect 37123 -2224 37187 -2160
rect 45110 -2224 45174 -2160
rect 10259 -2468 10323 -2404
rect 16406 -2468 16470 -2404
rect 17267 -2468 17331 -2404
rect 23894 -2468 23958 -2404
rect 27779 -2468 27843 -2404
rect 35126 -2468 35190 -2404
rect 35955 -2468 36019 -2404
rect 43862 -2468 43926 -2404
rect 6755 -2712 6819 -2648
rect 43577 -2712 43641 -2648
rect 44131 -2712 44195 -2648
rect 52598 -2712 52662 -2648
rect 4419 -2956 4483 -2892
rect 23609 -2956 23673 -2892
rect 26611 -2956 26675 -2892
rect 33878 -2956 33942 -2892
rect 34787 -2956 34851 -2892
rect 42614 -2956 42678 -2892
rect 42963 -2956 43027 -2892
rect 51350 -2956 51414 -2892
rect 3251 -3897 3315 -3893
rect 3251 -3953 3255 -3897
rect 3255 -3953 3311 -3897
rect 3311 -3953 3315 -3897
rect 3251 -3957 3315 -3953
rect 4419 -3897 4483 -3893
rect 4419 -3953 4423 -3897
rect 4423 -3953 4479 -3897
rect 4479 -3953 4483 -3897
rect 4419 -3957 4483 -3953
rect 5587 -3897 5651 -3893
rect 5587 -3953 5591 -3897
rect 5591 -3953 5647 -3897
rect 5647 -3953 5651 -3897
rect 5587 -3957 5651 -3953
rect 6755 -3897 6819 -3893
rect 6755 -3953 6759 -3897
rect 6759 -3953 6815 -3897
rect 6815 -3953 6819 -3897
rect 6755 -3957 6819 -3953
rect 7923 -3897 7987 -3893
rect 7923 -3953 7927 -3897
rect 7927 -3953 7983 -3897
rect 7983 -3953 7987 -3897
rect 7923 -3957 7987 -3953
rect 9091 -3897 9155 -3893
rect 9091 -3953 9095 -3897
rect 9095 -3953 9151 -3897
rect 9151 -3953 9155 -3897
rect 9091 -3957 9155 -3953
rect 10259 -3897 10323 -3893
rect 10259 -3953 10263 -3897
rect 10263 -3953 10319 -3897
rect 10319 -3953 10323 -3897
rect 10259 -3957 10323 -3953
rect 11427 -3897 11491 -3893
rect 11427 -3953 11431 -3897
rect 11431 -3953 11487 -3897
rect 11487 -3953 11491 -3897
rect 11427 -3957 11491 -3953
rect 12595 -3897 12659 -3893
rect 12595 -3953 12599 -3897
rect 12599 -3953 12655 -3897
rect 12655 -3953 12659 -3897
rect 12595 -3957 12659 -3953
rect 13763 -3897 13827 -3893
rect 13763 -3953 13767 -3897
rect 13767 -3953 13823 -3897
rect 13823 -3953 13827 -3897
rect 13763 -3957 13827 -3953
rect 14931 -3897 14995 -3893
rect 14931 -3953 14935 -3897
rect 14935 -3953 14991 -3897
rect 14991 -3953 14995 -3897
rect 14931 -3957 14995 -3953
rect 16099 -3897 16163 -3893
rect 16099 -3953 16103 -3897
rect 16103 -3953 16159 -3897
rect 16159 -3953 16163 -3897
rect 16099 -3957 16163 -3953
rect 17267 -3897 17331 -3893
rect 17267 -3953 17271 -3897
rect 17271 -3953 17327 -3897
rect 17327 -3953 17331 -3897
rect 17267 -3957 17331 -3953
rect 18435 -3897 18499 -3893
rect 18435 -3953 18439 -3897
rect 18439 -3953 18495 -3897
rect 18495 -3953 18499 -3897
rect 18435 -3957 18499 -3953
rect 19603 -3897 19667 -3893
rect 19603 -3953 19607 -3897
rect 19607 -3953 19663 -3897
rect 19663 -3953 19667 -3897
rect 19603 -3957 19667 -3953
rect 20771 -3897 20835 -3893
rect 20771 -3953 20775 -3897
rect 20775 -3953 20831 -3897
rect 20831 -3953 20835 -3897
rect 20771 -3957 20835 -3953
rect 21939 -3897 22003 -3893
rect 21939 -3953 21943 -3897
rect 21943 -3953 21999 -3897
rect 21999 -3953 22003 -3897
rect 21939 -3957 22003 -3953
rect 23107 -3897 23171 -3893
rect 23107 -3953 23111 -3897
rect 23111 -3953 23167 -3897
rect 23167 -3953 23171 -3897
rect 23107 -3957 23171 -3953
rect 24275 -3897 24339 -3893
rect 24275 -3953 24279 -3897
rect 24279 -3953 24335 -3897
rect 24335 -3953 24339 -3897
rect 24275 -3957 24339 -3953
rect 25443 -3897 25507 -3893
rect 25443 -3953 25447 -3897
rect 25447 -3953 25503 -3897
rect 25503 -3953 25507 -3897
rect 25443 -3957 25507 -3953
rect 26611 -3897 26675 -3893
rect 26611 -3953 26615 -3897
rect 26615 -3953 26671 -3897
rect 26671 -3953 26675 -3897
rect 26611 -3957 26675 -3953
rect 27779 -3897 27843 -3893
rect 27779 -3953 27783 -3897
rect 27783 -3953 27839 -3897
rect 27839 -3953 27843 -3897
rect 27779 -3957 27843 -3953
rect 28947 -3897 29011 -3893
rect 28947 -3953 28951 -3897
rect 28951 -3953 29007 -3897
rect 29007 -3953 29011 -3897
rect 28947 -3957 29011 -3953
rect 30115 -3897 30179 -3893
rect 30115 -3953 30119 -3897
rect 30119 -3953 30175 -3897
rect 30175 -3953 30179 -3897
rect 30115 -3957 30179 -3953
rect 31283 -3897 31347 -3893
rect 31283 -3953 31287 -3897
rect 31287 -3953 31343 -3897
rect 31343 -3953 31347 -3897
rect 31283 -3957 31347 -3953
rect 32451 -3897 32515 -3893
rect 32451 -3953 32455 -3897
rect 32455 -3953 32511 -3897
rect 32511 -3953 32515 -3897
rect 32451 -3957 32515 -3953
rect 33619 -3897 33683 -3893
rect 33619 -3953 33623 -3897
rect 33623 -3953 33679 -3897
rect 33679 -3953 33683 -3897
rect 33619 -3957 33683 -3953
rect 34787 -3897 34851 -3893
rect 34787 -3953 34791 -3897
rect 34791 -3953 34847 -3897
rect 34847 -3953 34851 -3897
rect 34787 -3957 34851 -3953
rect 35955 -3897 36019 -3893
rect 35955 -3953 35959 -3897
rect 35959 -3953 36015 -3897
rect 36015 -3953 36019 -3897
rect 35955 -3957 36019 -3953
rect 37123 -3897 37187 -3893
rect 37123 -3953 37127 -3897
rect 37127 -3953 37183 -3897
rect 37183 -3953 37187 -3897
rect 37123 -3957 37187 -3953
rect 38291 -3897 38355 -3893
rect 38291 -3953 38295 -3897
rect 38295 -3953 38351 -3897
rect 38351 -3953 38355 -3897
rect 38291 -3957 38355 -3953
rect 39459 -3897 39523 -3893
rect 39459 -3953 39463 -3897
rect 39463 -3953 39519 -3897
rect 39519 -3953 39523 -3897
rect 39459 -3957 39523 -3953
rect 40627 -3897 40691 -3893
rect 40627 -3953 40631 -3897
rect 40631 -3953 40687 -3897
rect 40687 -3953 40691 -3897
rect 40627 -3957 40691 -3953
rect 41795 -3897 41859 -3893
rect 41795 -3953 41799 -3897
rect 41799 -3953 41855 -3897
rect 41855 -3953 41859 -3897
rect 41795 -3957 41859 -3953
rect 42963 -3897 43027 -3893
rect 42963 -3953 42967 -3897
rect 42967 -3953 43023 -3897
rect 43023 -3953 43027 -3897
rect 42963 -3957 43027 -3953
rect 44131 -3897 44195 -3893
rect 44131 -3953 44135 -3897
rect 44135 -3953 44191 -3897
rect 44191 -3953 44195 -3897
rect 44131 -3957 44195 -3953
<< metal4 >>
rect 13909 1457 13975 1458
rect 13909 1393 13910 1457
rect 13974 1393 13975 1457
rect 13909 1392 13975 1393
rect 15157 1457 15223 1458
rect 15157 1393 15158 1457
rect 15222 1393 15223 1457
rect 15157 1392 15223 1393
rect 16405 1457 16471 1458
rect 16405 1393 16406 1457
rect 16470 1393 16471 1457
rect 16405 1392 16471 1393
rect 17653 1457 17719 1458
rect 17653 1393 17654 1457
rect 17718 1393 17719 1457
rect 17653 1392 17719 1393
rect 18901 1457 18967 1458
rect 18901 1393 18902 1457
rect 18966 1393 18967 1457
rect 18901 1392 18967 1393
rect 20149 1457 20215 1458
rect 20149 1393 20150 1457
rect 20214 1393 20215 1457
rect 20149 1392 20215 1393
rect 21397 1457 21463 1458
rect 21397 1393 21398 1457
rect 21462 1393 21463 1457
rect 21397 1392 21463 1393
rect 22645 1457 22711 1458
rect 22645 1393 22646 1457
rect 22710 1393 22711 1457
rect 22645 1392 22711 1393
rect 23893 1457 23959 1458
rect 23893 1393 23894 1457
rect 23958 1393 23959 1457
rect 23893 1392 23959 1393
rect 25141 1457 25207 1458
rect 25141 1393 25142 1457
rect 25206 1393 25207 1457
rect 25141 1392 25207 1393
rect 26389 1457 26455 1458
rect 26389 1393 26390 1457
rect 26454 1393 26455 1457
rect 26389 1392 26455 1393
rect 27637 1457 27703 1458
rect 27637 1393 27638 1457
rect 27702 1393 27703 1457
rect 27637 1392 27703 1393
rect 28885 1457 28951 1458
rect 28885 1393 28886 1457
rect 28950 1393 28951 1457
rect 28885 1392 28951 1393
rect 30133 1457 30199 1458
rect 30133 1393 30134 1457
rect 30198 1393 30199 1457
rect 30133 1392 30199 1393
rect 31381 1457 31447 1458
rect 31381 1393 31382 1457
rect 31446 1393 31447 1457
rect 31381 1392 31447 1393
rect 32629 1457 32695 1458
rect 32629 1393 32630 1457
rect 32694 1393 32695 1457
rect 32629 1392 32695 1393
rect 33877 1457 33943 1458
rect 33877 1393 33878 1457
rect 33942 1393 33943 1457
rect 33877 1392 33943 1393
rect 35125 1457 35191 1458
rect 35125 1393 35126 1457
rect 35190 1393 35191 1457
rect 35125 1392 35191 1393
rect 36373 1457 36439 1458
rect 36373 1393 36374 1457
rect 36438 1393 36439 1457
rect 36373 1392 36439 1393
rect 37621 1457 37687 1458
rect 37621 1393 37622 1457
rect 37686 1393 37687 1457
rect 37621 1392 37687 1393
rect 38869 1457 38935 1458
rect 38869 1393 38870 1457
rect 38934 1393 38935 1457
rect 38869 1392 38935 1393
rect 40117 1457 40183 1458
rect 40117 1393 40118 1457
rect 40182 1393 40183 1457
rect 40117 1392 40183 1393
rect 41365 1457 41431 1458
rect 41365 1393 41366 1457
rect 41430 1393 41431 1457
rect 41365 1392 41431 1393
rect 42613 1457 42679 1458
rect 42613 1393 42614 1457
rect 42678 1393 42679 1457
rect 42613 1392 42679 1393
rect 43861 1457 43927 1458
rect 43861 1393 43862 1457
rect 43926 1393 43927 1457
rect 43861 1392 43927 1393
rect 45109 1457 45175 1458
rect 45109 1393 45110 1457
rect 45174 1393 45175 1457
rect 45109 1392 45175 1393
rect 46357 1457 46423 1458
rect 46357 1393 46358 1457
rect 46422 1393 46423 1457
rect 46357 1392 46423 1393
rect 47605 1457 47671 1458
rect 47605 1393 47606 1457
rect 47670 1393 47671 1457
rect 47605 1392 47671 1393
rect 48853 1457 48919 1458
rect 48853 1393 48854 1457
rect 48918 1393 48919 1457
rect 48853 1392 48919 1393
rect 50101 1457 50167 1458
rect 50101 1393 50102 1457
rect 50166 1393 50167 1457
rect 50101 1392 50167 1393
rect 51349 1457 51415 1458
rect 51349 1393 51350 1457
rect 51414 1393 51415 1457
rect 51349 1392 51415 1393
rect 52597 1457 52663 1458
rect 52597 1393 52598 1457
rect 52662 1393 52663 1457
rect 52597 1392 52663 1393
rect 13624 337 13690 338
rect 13624 273 13625 337
rect 13689 273 13690 337
rect 13624 272 13690 273
rect 9090 -696 9156 -695
rect 9090 -760 9091 -696
rect 9155 -760 9156 -696
rect 9090 -761 9156 -760
rect 5586 -940 5652 -939
rect 5586 -1004 5587 -940
rect 5651 -1004 5652 -940
rect 5586 -1005 5652 -1004
rect 3250 -1428 3316 -1427
rect 3250 -1492 3251 -1428
rect 3315 -1492 3316 -1428
rect 3250 -1493 3316 -1492
rect 3253 -3892 3313 -1493
rect 4418 -2892 4484 -2891
rect 4418 -2956 4419 -2892
rect 4483 -2956 4484 -2892
rect 4418 -2957 4484 -2956
rect 4421 -3892 4481 -2957
rect 5589 -3892 5649 -1005
rect 7922 -1184 7988 -1183
rect 7922 -1248 7923 -1184
rect 7987 -1248 7988 -1184
rect 7922 -1249 7988 -1248
rect 6754 -2648 6820 -2647
rect 6754 -2712 6755 -2648
rect 6819 -2712 6820 -2648
rect 6754 -2713 6820 -2712
rect 6757 -3892 6817 -2713
rect 7925 -3892 7985 -1249
rect 9093 -3892 9153 -761
rect 13627 -1427 13687 272
rect 13912 -1183 13972 1392
rect 15160 -695 15220 1392
rect 15157 -696 15223 -695
rect 15157 -760 15158 -696
rect 15222 -760 15223 -696
rect 15157 -761 15223 -760
rect 13909 -1184 13975 -1183
rect 13909 -1248 13910 -1184
rect 13974 -1248 13975 -1184
rect 13909 -1249 13975 -1248
rect 16098 -1184 16164 -1183
rect 16098 -1248 16099 -1184
rect 16163 -1248 16164 -1184
rect 16098 -1249 16164 -1248
rect 13624 -1428 13690 -1427
rect 13624 -1492 13625 -1428
rect 13689 -1492 13690 -1428
rect 13624 -1493 13690 -1492
rect 14930 -1428 14996 -1427
rect 14930 -1492 14931 -1428
rect 14995 -1492 14996 -1428
rect 14930 -1493 14996 -1492
rect 13762 -1672 13828 -1671
rect 13762 -1736 13763 -1672
rect 13827 -1736 13828 -1672
rect 13762 -1737 13828 -1736
rect 12594 -1916 12660 -1915
rect 12594 -1980 12595 -1916
rect 12659 -1980 12660 -1916
rect 12594 -1981 12660 -1980
rect 11426 -2160 11492 -2159
rect 11426 -2224 11427 -2160
rect 11491 -2224 11492 -2160
rect 11426 -2225 11492 -2224
rect 10258 -2404 10324 -2403
rect 10258 -2468 10259 -2404
rect 10323 -2468 10324 -2404
rect 10258 -2469 10324 -2468
rect 10261 -3892 10321 -2469
rect 11429 -3892 11489 -2225
rect 12597 -3892 12657 -1981
rect 13765 -3892 13825 -1737
rect 14933 -3892 14993 -1493
rect 16101 -3892 16161 -1249
rect 16408 -2403 16468 1392
rect 17656 -2159 17716 1392
rect 18904 -1915 18964 1392
rect 20152 -1671 20212 1392
rect 21400 -1427 21460 1392
rect 22648 -1183 22708 1392
rect 23608 337 23674 338
rect 23608 273 23609 337
rect 23673 273 23674 337
rect 23608 272 23674 273
rect 22645 -1184 22711 -1183
rect 22645 -1248 22646 -1184
rect 22710 -1248 22711 -1184
rect 22645 -1249 22711 -1248
rect 23106 -1184 23172 -1183
rect 23106 -1248 23107 -1184
rect 23171 -1248 23172 -1184
rect 23106 -1249 23172 -1248
rect 21397 -1428 21463 -1427
rect 21397 -1492 21398 -1428
rect 21462 -1492 21463 -1428
rect 21397 -1493 21463 -1492
rect 21938 -1428 22004 -1427
rect 21938 -1492 21939 -1428
rect 22003 -1492 22004 -1428
rect 21938 -1493 22004 -1492
rect 20149 -1672 20215 -1671
rect 20149 -1736 20150 -1672
rect 20214 -1736 20215 -1672
rect 20149 -1737 20215 -1736
rect 20770 -1672 20836 -1671
rect 20770 -1736 20771 -1672
rect 20835 -1736 20836 -1672
rect 20770 -1737 20836 -1736
rect 18901 -1916 18967 -1915
rect 18901 -1980 18902 -1916
rect 18966 -1980 18967 -1916
rect 18901 -1981 18967 -1980
rect 19602 -1916 19668 -1915
rect 19602 -1980 19603 -1916
rect 19667 -1980 19668 -1916
rect 19602 -1981 19668 -1980
rect 17653 -2160 17719 -2159
rect 17653 -2224 17654 -2160
rect 17718 -2224 17719 -2160
rect 17653 -2225 17719 -2224
rect 18434 -2160 18500 -2159
rect 18434 -2224 18435 -2160
rect 18499 -2224 18500 -2160
rect 18434 -2225 18500 -2224
rect 16405 -2404 16471 -2403
rect 16405 -2468 16406 -2404
rect 16470 -2468 16471 -2404
rect 16405 -2469 16471 -2468
rect 17266 -2404 17332 -2403
rect 17266 -2468 17267 -2404
rect 17331 -2468 17332 -2404
rect 17266 -2469 17332 -2468
rect 17269 -3892 17329 -2469
rect 18437 -3892 18497 -2225
rect 19605 -3892 19665 -1981
rect 20773 -3892 20833 -1737
rect 21941 -3892 22001 -1493
rect 23109 -3892 23169 -1249
rect 23611 -2891 23671 272
rect 23896 -2403 23956 1392
rect 24274 -696 24340 -695
rect 24274 -760 24275 -696
rect 24339 -760 24340 -696
rect 24274 -761 24340 -760
rect 23893 -2404 23959 -2403
rect 23893 -2468 23894 -2404
rect 23958 -2468 23959 -2404
rect 23893 -2469 23959 -2468
rect 23608 -2892 23674 -2891
rect 23608 -2956 23609 -2892
rect 23673 -2956 23674 -2892
rect 23608 -2957 23674 -2956
rect 24277 -3892 24337 -761
rect 25144 -2159 25204 1392
rect 25442 -452 25508 -451
rect 25442 -516 25443 -452
rect 25507 -516 25508 -452
rect 25442 -517 25508 -516
rect 25141 -2160 25207 -2159
rect 25141 -2224 25142 -2160
rect 25206 -2224 25207 -2160
rect 25141 -2225 25207 -2224
rect 25445 -3892 25505 -517
rect 26392 -1915 26452 1392
rect 27640 -1671 27700 1392
rect 28888 -1427 28948 1392
rect 30136 -1183 30196 1392
rect 31384 -695 31444 1392
rect 32632 -451 32692 1392
rect 33592 337 33658 338
rect 33592 273 33593 337
rect 33657 273 33658 337
rect 33592 272 33658 273
rect 32629 -452 32695 -451
rect 32629 -516 32630 -452
rect 32694 -516 32695 -452
rect 32629 -517 32695 -516
rect 31381 -696 31447 -695
rect 31381 -760 31382 -696
rect 31446 -760 31447 -696
rect 31381 -761 31447 -760
rect 33595 -939 33655 272
rect 33592 -940 33658 -939
rect 33592 -1004 33593 -940
rect 33657 -1004 33658 -940
rect 33592 -1005 33658 -1004
rect 30133 -1184 30199 -1183
rect 30133 -1248 30134 -1184
rect 30198 -1248 30199 -1184
rect 30133 -1249 30199 -1248
rect 33618 -1184 33684 -1183
rect 33618 -1248 33619 -1184
rect 33683 -1248 33684 -1184
rect 33618 -1249 33684 -1248
rect 28885 -1428 28951 -1427
rect 28885 -1492 28886 -1428
rect 28950 -1492 28951 -1428
rect 28885 -1493 28951 -1492
rect 32450 -1428 32516 -1427
rect 32450 -1492 32451 -1428
rect 32515 -1492 32516 -1428
rect 32450 -1493 32516 -1492
rect 27637 -1672 27703 -1671
rect 27637 -1736 27638 -1672
rect 27702 -1736 27703 -1672
rect 27637 -1737 27703 -1736
rect 31282 -1672 31348 -1671
rect 31282 -1736 31283 -1672
rect 31347 -1736 31348 -1672
rect 31282 -1737 31348 -1736
rect 26389 -1916 26455 -1915
rect 26389 -1980 26390 -1916
rect 26454 -1980 26455 -1916
rect 26389 -1981 26455 -1980
rect 30114 -1916 30180 -1915
rect 30114 -1980 30115 -1916
rect 30179 -1980 30180 -1916
rect 30114 -1981 30180 -1980
rect 28946 -2160 29012 -2159
rect 28946 -2224 28947 -2160
rect 29011 -2224 29012 -2160
rect 28946 -2225 29012 -2224
rect 27778 -2404 27844 -2403
rect 27778 -2468 27779 -2404
rect 27843 -2468 27844 -2404
rect 27778 -2469 27844 -2468
rect 26610 -2892 26676 -2891
rect 26610 -2956 26611 -2892
rect 26675 -2956 26676 -2892
rect 26610 -2957 26676 -2956
rect 26613 -3892 26673 -2957
rect 27781 -3892 27841 -2469
rect 28949 -3892 29009 -2225
rect 30117 -3892 30177 -1981
rect 31285 -3892 31345 -1737
rect 32453 -3892 32513 -1493
rect 33621 -3892 33681 -1249
rect 33880 -2891 33940 1392
rect 35128 -2403 35188 1392
rect 36376 -2159 36436 1392
rect 37624 -1915 37684 1392
rect 38872 -1671 38932 1392
rect 40120 -1427 40180 1392
rect 41368 -1183 41428 1392
rect 41365 -1184 41431 -1183
rect 41365 -1248 41366 -1184
rect 41430 -1248 41431 -1184
rect 41365 -1249 41431 -1248
rect 41794 -1184 41860 -1183
rect 41794 -1248 41795 -1184
rect 41859 -1248 41860 -1184
rect 41794 -1249 41860 -1248
rect 40117 -1428 40183 -1427
rect 40117 -1492 40118 -1428
rect 40182 -1492 40183 -1428
rect 40117 -1493 40183 -1492
rect 40626 -1428 40692 -1427
rect 40626 -1492 40627 -1428
rect 40691 -1492 40692 -1428
rect 40626 -1493 40692 -1492
rect 38869 -1672 38935 -1671
rect 38869 -1736 38870 -1672
rect 38934 -1736 38935 -1672
rect 38869 -1737 38935 -1736
rect 39458 -1672 39524 -1671
rect 39458 -1736 39459 -1672
rect 39523 -1736 39524 -1672
rect 39458 -1737 39524 -1736
rect 37621 -1916 37687 -1915
rect 37621 -1980 37622 -1916
rect 37686 -1980 37687 -1916
rect 37621 -1981 37687 -1980
rect 38290 -1916 38356 -1915
rect 38290 -1980 38291 -1916
rect 38355 -1980 38356 -1916
rect 38290 -1981 38356 -1980
rect 36373 -2160 36439 -2159
rect 36373 -2224 36374 -2160
rect 36438 -2224 36439 -2160
rect 36373 -2225 36439 -2224
rect 37122 -2160 37188 -2159
rect 37122 -2224 37123 -2160
rect 37187 -2224 37188 -2160
rect 37122 -2225 37188 -2224
rect 35125 -2404 35191 -2403
rect 35125 -2468 35126 -2404
rect 35190 -2468 35191 -2404
rect 35125 -2469 35191 -2468
rect 35954 -2404 36020 -2403
rect 35954 -2468 35955 -2404
rect 36019 -2468 36020 -2404
rect 35954 -2469 36020 -2468
rect 33877 -2892 33943 -2891
rect 33877 -2956 33878 -2892
rect 33942 -2956 33943 -2892
rect 33877 -2957 33943 -2956
rect 34786 -2892 34852 -2891
rect 34786 -2956 34787 -2892
rect 34851 -2956 34852 -2892
rect 34786 -2957 34852 -2956
rect 34789 -3892 34849 -2957
rect 35957 -3892 36017 -2469
rect 37125 -3892 37185 -2225
rect 38293 -3892 38353 -1981
rect 39461 -3892 39521 -1737
rect 40629 -3892 40689 -1493
rect 41797 -3892 41857 -1249
rect 42616 -2891 42676 1392
rect 43576 337 43642 338
rect 43576 273 43577 337
rect 43641 273 43642 337
rect 43576 272 43642 273
rect 43579 -2647 43639 272
rect 43864 -2403 43924 1392
rect 45112 -2159 45172 1392
rect 46360 -1915 46420 1392
rect 47608 -1671 47668 1392
rect 48856 -1427 48916 1392
rect 50104 -1183 50164 1392
rect 50101 -1184 50167 -1183
rect 50101 -1248 50102 -1184
rect 50166 -1248 50167 -1184
rect 50101 -1249 50167 -1248
rect 48853 -1428 48919 -1427
rect 48853 -1492 48854 -1428
rect 48918 -1492 48919 -1428
rect 48853 -1493 48919 -1492
rect 47605 -1672 47671 -1671
rect 47605 -1736 47606 -1672
rect 47670 -1736 47671 -1672
rect 47605 -1737 47671 -1736
rect 46357 -1916 46423 -1915
rect 46357 -1980 46358 -1916
rect 46422 -1980 46423 -1916
rect 46357 -1981 46423 -1980
rect 45109 -2160 45175 -2159
rect 45109 -2224 45110 -2160
rect 45174 -2224 45175 -2160
rect 45109 -2225 45175 -2224
rect 43861 -2404 43927 -2403
rect 43861 -2468 43862 -2404
rect 43926 -2468 43927 -2404
rect 43861 -2469 43927 -2468
rect 43576 -2648 43642 -2647
rect 43576 -2712 43577 -2648
rect 43641 -2712 43642 -2648
rect 43576 -2713 43642 -2712
rect 44130 -2648 44196 -2647
rect 44130 -2712 44131 -2648
rect 44195 -2712 44196 -2648
rect 44130 -2713 44196 -2712
rect 42613 -2892 42679 -2891
rect 42613 -2956 42614 -2892
rect 42678 -2956 42679 -2892
rect 42613 -2957 42679 -2956
rect 42962 -2892 43028 -2891
rect 42962 -2956 42963 -2892
rect 43027 -2956 43028 -2892
rect 42962 -2957 43028 -2956
rect 42965 -3892 43025 -2957
rect 44133 -3892 44193 -2713
rect 51352 -2891 51412 1392
rect 52600 -2647 52660 1392
rect 52597 -2648 52663 -2647
rect 52597 -2712 52598 -2648
rect 52662 -2712 52663 -2648
rect 52597 -2713 52663 -2712
rect 51349 -2892 51415 -2891
rect 51349 -2956 51350 -2892
rect 51414 -2956 51415 -2892
rect 51349 -2957 51415 -2956
rect 3250 -3893 3316 -3892
rect 3250 -3957 3251 -3893
rect 3315 -3957 3316 -3893
rect 3250 -3958 3316 -3957
rect 4418 -3893 4484 -3892
rect 4418 -3957 4419 -3893
rect 4483 -3957 4484 -3893
rect 4418 -3958 4484 -3957
rect 5586 -3893 5652 -3892
rect 5586 -3957 5587 -3893
rect 5651 -3957 5652 -3893
rect 5586 -3958 5652 -3957
rect 6754 -3893 6820 -3892
rect 6754 -3957 6755 -3893
rect 6819 -3957 6820 -3893
rect 6754 -3958 6820 -3957
rect 7922 -3893 7988 -3892
rect 7922 -3957 7923 -3893
rect 7987 -3957 7988 -3893
rect 7922 -3958 7988 -3957
rect 9090 -3893 9156 -3892
rect 9090 -3957 9091 -3893
rect 9155 -3957 9156 -3893
rect 9090 -3958 9156 -3957
rect 10258 -3893 10324 -3892
rect 10258 -3957 10259 -3893
rect 10323 -3957 10324 -3893
rect 10258 -3958 10324 -3957
rect 11426 -3893 11492 -3892
rect 11426 -3957 11427 -3893
rect 11491 -3957 11492 -3893
rect 11426 -3958 11492 -3957
rect 12594 -3893 12660 -3892
rect 12594 -3957 12595 -3893
rect 12659 -3957 12660 -3893
rect 12594 -3958 12660 -3957
rect 13762 -3893 13828 -3892
rect 13762 -3957 13763 -3893
rect 13827 -3957 13828 -3893
rect 13762 -3958 13828 -3957
rect 14930 -3893 14996 -3892
rect 14930 -3957 14931 -3893
rect 14995 -3957 14996 -3893
rect 14930 -3958 14996 -3957
rect 16098 -3893 16164 -3892
rect 16098 -3957 16099 -3893
rect 16163 -3957 16164 -3893
rect 16098 -3958 16164 -3957
rect 17266 -3893 17332 -3892
rect 17266 -3957 17267 -3893
rect 17331 -3957 17332 -3893
rect 17266 -3958 17332 -3957
rect 18434 -3893 18500 -3892
rect 18434 -3957 18435 -3893
rect 18499 -3957 18500 -3893
rect 18434 -3958 18500 -3957
rect 19602 -3893 19668 -3892
rect 19602 -3957 19603 -3893
rect 19667 -3957 19668 -3893
rect 19602 -3958 19668 -3957
rect 20770 -3893 20836 -3892
rect 20770 -3957 20771 -3893
rect 20835 -3957 20836 -3893
rect 20770 -3958 20836 -3957
rect 21938 -3893 22004 -3892
rect 21938 -3957 21939 -3893
rect 22003 -3957 22004 -3893
rect 21938 -3958 22004 -3957
rect 23106 -3893 23172 -3892
rect 23106 -3957 23107 -3893
rect 23171 -3957 23172 -3893
rect 23106 -3958 23172 -3957
rect 24274 -3893 24340 -3892
rect 24274 -3957 24275 -3893
rect 24339 -3957 24340 -3893
rect 24274 -3958 24340 -3957
rect 25442 -3893 25508 -3892
rect 25442 -3957 25443 -3893
rect 25507 -3957 25508 -3893
rect 25442 -3958 25508 -3957
rect 26610 -3893 26676 -3892
rect 26610 -3957 26611 -3893
rect 26675 -3957 26676 -3893
rect 26610 -3958 26676 -3957
rect 27778 -3893 27844 -3892
rect 27778 -3957 27779 -3893
rect 27843 -3957 27844 -3893
rect 27778 -3958 27844 -3957
rect 28946 -3893 29012 -3892
rect 28946 -3957 28947 -3893
rect 29011 -3957 29012 -3893
rect 28946 -3958 29012 -3957
rect 30114 -3893 30180 -3892
rect 30114 -3957 30115 -3893
rect 30179 -3957 30180 -3893
rect 30114 -3958 30180 -3957
rect 31282 -3893 31348 -3892
rect 31282 -3957 31283 -3893
rect 31347 -3957 31348 -3893
rect 31282 -3958 31348 -3957
rect 32450 -3893 32516 -3892
rect 32450 -3957 32451 -3893
rect 32515 -3957 32516 -3893
rect 32450 -3958 32516 -3957
rect 33618 -3893 33684 -3892
rect 33618 -3957 33619 -3893
rect 33683 -3957 33684 -3893
rect 33618 -3958 33684 -3957
rect 34786 -3893 34852 -3892
rect 34786 -3957 34787 -3893
rect 34851 -3957 34852 -3893
rect 34786 -3958 34852 -3957
rect 35954 -3893 36020 -3892
rect 35954 -3957 35955 -3893
rect 36019 -3957 36020 -3893
rect 35954 -3958 36020 -3957
rect 37122 -3893 37188 -3892
rect 37122 -3957 37123 -3893
rect 37187 -3957 37188 -3893
rect 37122 -3958 37188 -3957
rect 38290 -3893 38356 -3892
rect 38290 -3957 38291 -3893
rect 38355 -3957 38356 -3893
rect 38290 -3958 38356 -3957
rect 39458 -3893 39524 -3892
rect 39458 -3957 39459 -3893
rect 39523 -3957 39524 -3893
rect 39458 -3958 39524 -3957
rect 40626 -3893 40692 -3892
rect 40626 -3957 40627 -3893
rect 40691 -3957 40692 -3893
rect 40626 -3958 40692 -3957
rect 41794 -3893 41860 -3892
rect 41794 -3957 41795 -3893
rect 41859 -3957 41860 -3893
rect 41794 -3958 41860 -3957
rect 42962 -3893 43028 -3892
rect 42962 -3957 42963 -3893
rect 43027 -3957 43028 -3893
rect 42962 -3958 43028 -3957
rect 44130 -3893 44196 -3892
rect 44130 -3957 44131 -3893
rect 44195 -3957 44196 -3893
rect 44130 -3958 44196 -3957
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_0
timestamp 1666464484
transform 1 0 12594 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_1
timestamp 1666464484
transform 1 0 3250 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_2
timestamp 1666464484
transform 1 0 13624 0 1 268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_3
timestamp 1666464484
transform 1 0 4418 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_4
timestamp 1666464484
transform 1 0 9090 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_5
timestamp 1666464484
transform 1 0 15157 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_6
timestamp 1666464484
transform 1 0 5586 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_7
timestamp 1666464484
transform 1 0 7922 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_8
timestamp 1666464484
transform 1 0 13909 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_9
timestamp 1666464484
transform 1 0 6754 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_10
timestamp 1666464484
transform 1 0 11426 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_11
timestamp 1666464484
transform 1 0 14930 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_12
timestamp 1666464484
transform 1 0 13762 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_13
timestamp 1666464484
transform 1 0 10258 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_14
timestamp 1666464484
transform 1 0 25442 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_15
timestamp 1666464484
transform 1 0 20149 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_16
timestamp 1666464484
transform 1 0 24274 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_17
timestamp 1666464484
transform 1 0 23608 0 1 268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_18
timestamp 1666464484
transform 1 0 27778 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_19
timestamp 1666464484
transform 1 0 26610 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_20
timestamp 1666464484
transform 1 0 19602 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_21
timestamp 1666464484
transform 1 0 26389 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_22
timestamp 1666464484
transform 1 0 23106 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_23
timestamp 1666464484
transform 1 0 16098 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_24
timestamp 1666464484
transform 1 0 22645 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_25
timestamp 1666464484
transform 1 0 18901 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_26
timestamp 1666464484
transform 1 0 17266 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_27
timestamp 1666464484
transform 1 0 23893 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_28
timestamp 1666464484
transform 1 0 16405 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_29
timestamp 1666464484
transform 1 0 21938 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_30
timestamp 1666464484
transform 1 0 21397 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_31
timestamp 1666464484
transform 1 0 18434 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_32
timestamp 1666464484
transform 1 0 25141 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_33
timestamp 1666464484
transform 1 0 17653 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_34
timestamp 1666464484
transform 1 0 20770 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_35
timestamp 1666464484
transform 1 0 27637 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_36
timestamp 1666464484
transform 1 0 32629 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_37
timestamp 1666464484
transform 1 0 31381 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_38
timestamp 1666464484
transform 1 0 33592 0 1 268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_39
timestamp 1666464484
transform 1 0 37122 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_40
timestamp 1666464484
transform 1 0 33877 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_41
timestamp 1666464484
transform 1 0 33618 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_42
timestamp 1666464484
transform 1 0 28946 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_43
timestamp 1666464484
transform 1 0 30133 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_44
timestamp 1666464484
transform 1 0 36373 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_45
timestamp 1666464484
transform 1 0 35954 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_46
timestamp 1666464484
transform 1 0 32450 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_47
timestamp 1666464484
transform 1 0 40117 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_48
timestamp 1666464484
transform 1 0 28885 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_49
timestamp 1666464484
transform 1 0 39458 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_50
timestamp 1666464484
transform 1 0 34786 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_51
timestamp 1666464484
transform 1 0 31282 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_52
timestamp 1666464484
transform 1 0 38869 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_53
timestamp 1666464484
transform 1 0 38290 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_54
timestamp 1666464484
transform 1 0 35125 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_55
timestamp 1666464484
transform 1 0 30114 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_56
timestamp 1666464484
transform 1 0 37621 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_57
timestamp 1666464484
transform 1 0 41794 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_58
timestamp 1666464484
transform 1 0 50101 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_59
timestamp 1666464484
transform 1 0 41365 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_60
timestamp 1666464484
transform 1 0 40626 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_61
timestamp 1666464484
transform 1 0 48853 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_62
timestamp 1666464484
transform 1 0 47605 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_63
timestamp 1666464484
transform 1 0 46357 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_64
timestamp 1666464484
transform 1 0 45109 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_65
timestamp 1666464484
transform 1 0 43861 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_66
timestamp 1666464484
transform 1 0 44130 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_67
timestamp 1666464484
transform 1 0 52597 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_68
timestamp 1666464484
transform 1 0 43576 0 1 268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_69
timestamp 1666464484
transform 1 0 42962 0 1 -3962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_70
timestamp 1666464484
transform 1 0 51349 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_71
timestamp 1666464484
transform 1 0 42613 0 1 1388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1666464484
transform 1 0 15158 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1666464484
transform 1 0 13910 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1666464484
transform 1 0 20150 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_3
timestamp 1666464484
transform 1 0 26390 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_4
timestamp 1666464484
transform 1 0 22646 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_5
timestamp 1666464484
transform 1 0 18902 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_6
timestamp 1666464484
transform 1 0 23894 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_7
timestamp 1666464484
transform 1 0 16406 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_8
timestamp 1666464484
transform 1 0 21398 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_9
timestamp 1666464484
transform 1 0 25142 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_10
timestamp 1666464484
transform 1 0 17654 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_11
timestamp 1666464484
transform 1 0 27638 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_12
timestamp 1666464484
transform 1 0 32630 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_13
timestamp 1666464484
transform 1 0 31382 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_14
timestamp 1666464484
transform 1 0 37622 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_15
timestamp 1666464484
transform 1 0 33878 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_16
timestamp 1666464484
transform 1 0 30134 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_17
timestamp 1666464484
transform 1 0 36374 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_18
timestamp 1666464484
transform 1 0 40118 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_19
timestamp 1666464484
transform 1 0 28886 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_20
timestamp 1666464484
transform 1 0 38870 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_21
timestamp 1666464484
transform 1 0 35126 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_22
timestamp 1666464484
transform 1 0 50102 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_23
timestamp 1666464484
transform 1 0 41366 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_24
timestamp 1666464484
transform 1 0 48854 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_25
timestamp 1666464484
transform 1 0 47606 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_26
timestamp 1666464484
transform 1 0 46358 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_27
timestamp 1666464484
transform 1 0 45110 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_28
timestamp 1666464484
transform 1 0 43862 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_29
timestamp 1666464484
transform 1 0 52598 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_30
timestamp 1666464484
transform 1 0 51350 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_31
timestamp 1666464484
transform 1 0 42614 0 1 1393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_0
timestamp 1666464484
transform 1 0 12589 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1
timestamp 1666464484
transform 1 0 12589 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2
timestamp 1666464484
transform 1 0 10253 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_3
timestamp 1666464484
transform 1 0 3245 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_4
timestamp 1666464484
transform 1 0 3245 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_5
timestamp 1666464484
transform 1 0 13619 0 1 272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_6
timestamp 1666464484
transform 1 0 13619 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_7
timestamp 1666464484
transform 1 0 11421 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_8
timestamp 1666464484
transform 1 0 7917 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_9
timestamp 1666464484
transform 1 0 4413 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_10
timestamp 1666464484
transform 1 0 9085 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_11
timestamp 1666464484
transform 1 0 9085 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_12
timestamp 1666464484
transform 1 0 15152 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_13
timestamp 1666464484
transform 1 0 15152 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_14
timestamp 1666464484
transform 1 0 5581 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_15
timestamp 1666464484
transform 1 0 5581 0 1 -1005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_16
timestamp 1666464484
transform 1 0 6749 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_17
timestamp 1666464484
transform 1 0 7917 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_18
timestamp 1666464484
transform 1 0 13904 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_19
timestamp 1666464484
transform 1 0 6749 0 1 -2713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_20
timestamp 1666464484
transform 1 0 13904 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_21
timestamp 1666464484
transform 1 0 4413 0 1 -2957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_22
timestamp 1666464484
transform 1 0 14925 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_23
timestamp 1666464484
transform 1 0 14925 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_24
timestamp 1666464484
transform 1 0 11421 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_25
timestamp 1666464484
transform 1 0 13757 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_26
timestamp 1666464484
transform 1 0 13757 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_27
timestamp 1666464484
transform 1 0 10253 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_28
timestamp 1666464484
transform 1 0 25437 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_29
timestamp 1666464484
transform 1 0 25437 0 1 -517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_30
timestamp 1666464484
transform 1 0 20144 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_31
timestamp 1666464484
transform 1 0 20144 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_32
timestamp 1666464484
transform 1 0 24269 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_33
timestamp 1666464484
transform 1 0 24269 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_34
timestamp 1666464484
transform 1 0 23603 0 1 -2957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_35
timestamp 1666464484
transform 1 0 26605 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_36
timestamp 1666464484
transform 1 0 27773 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_37
timestamp 1666464484
transform 1 0 27773 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_38
timestamp 1666464484
transform 1 0 26605 0 1 -2957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_39
timestamp 1666464484
transform 1 0 17261 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_40
timestamp 1666464484
transform 1 0 19597 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_41
timestamp 1666464484
transform 1 0 19597 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_42
timestamp 1666464484
transform 1 0 26384 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_43
timestamp 1666464484
transform 1 0 26384 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_44
timestamp 1666464484
transform 1 0 23101 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_45
timestamp 1666464484
transform 1 0 23101 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_46
timestamp 1666464484
transform 1 0 18896 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_47
timestamp 1666464484
transform 1 0 16093 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_48
timestamp 1666464484
transform 1 0 16093 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_49
timestamp 1666464484
transform 1 0 22640 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_50
timestamp 1666464484
transform 1 0 22640 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_51
timestamp 1666464484
transform 1 0 18896 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_52
timestamp 1666464484
transform 1 0 17261 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_53
timestamp 1666464484
transform 1 0 23888 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_54
timestamp 1666464484
transform 1 0 23888 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_55
timestamp 1666464484
transform 1 0 16400 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_56
timestamp 1666464484
transform 1 0 21933 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_57
timestamp 1666464484
transform 1 0 21933 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_58
timestamp 1666464484
transform 1 0 16400 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_59
timestamp 1666464484
transform 1 0 18429 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_60
timestamp 1666464484
transform 1 0 21392 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_61
timestamp 1666464484
transform 1 0 21392 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_62
timestamp 1666464484
transform 1 0 18429 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_63
timestamp 1666464484
transform 1 0 25136 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_64
timestamp 1666464484
transform 1 0 25136 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_65
timestamp 1666464484
transform 1 0 17648 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_66
timestamp 1666464484
transform 1 0 17648 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_67
timestamp 1666464484
transform 1 0 23603 0 1 272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_68
timestamp 1666464484
transform 1 0 20765 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_69
timestamp 1666464484
transform 1 0 20765 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_70
timestamp 1666464484
transform 1 0 27632 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_71
timestamp 1666464484
transform 1 0 27632 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_72
timestamp 1666464484
transform 1 0 32624 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_73
timestamp 1666464484
transform 1 0 32624 0 1 -517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_74
timestamp 1666464484
transform 1 0 31376 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_75
timestamp 1666464484
transform 1 0 31376 0 1 -761
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_76
timestamp 1666464484
transform 1 0 33587 0 1 272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_77
timestamp 1666464484
transform 1 0 33587 0 1 -1005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_78
timestamp 1666464484
transform 1 0 37616 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_79
timestamp 1666464484
transform 1 0 37117 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_80
timestamp 1666464484
transform 1 0 37117 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_81
timestamp 1666464484
transform 1 0 35120 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_82
timestamp 1666464484
transform 1 0 33613 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_83
timestamp 1666464484
transform 1 0 33613 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_84
timestamp 1666464484
transform 1 0 33872 0 1 -2957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_85
timestamp 1666464484
transform 1 0 28941 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_86
timestamp 1666464484
transform 1 0 30128 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_87
timestamp 1666464484
transform 1 0 30128 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_88
timestamp 1666464484
transform 1 0 28941 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_89
timestamp 1666464484
transform 1 0 36368 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_90
timestamp 1666464484
transform 1 0 36368 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_91
timestamp 1666464484
transform 1 0 35949 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_92
timestamp 1666464484
transform 1 0 32445 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_93
timestamp 1666464484
transform 1 0 32445 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_94
timestamp 1666464484
transform 1 0 40112 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_95
timestamp 1666464484
transform 1 0 40112 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_96
timestamp 1666464484
transform 1 0 28880 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_97
timestamp 1666464484
transform 1 0 28880 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_98
timestamp 1666464484
transform 1 0 39453 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_99
timestamp 1666464484
transform 1 0 39453 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_100
timestamp 1666464484
transform 1 0 35949 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_101
timestamp 1666464484
transform 1 0 34781 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_102
timestamp 1666464484
transform 1 0 34781 0 1 -2957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_103
timestamp 1666464484
transform 1 0 31277 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_104
timestamp 1666464484
transform 1 0 31277 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_105
timestamp 1666464484
transform 1 0 38864 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_106
timestamp 1666464484
transform 1 0 38864 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_107
timestamp 1666464484
transform 1 0 38285 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_108
timestamp 1666464484
transform 1 0 38285 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_109
timestamp 1666464484
transform 1 0 33872 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_110
timestamp 1666464484
transform 1 0 35120 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_111
timestamp 1666464484
transform 1 0 30109 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_112
timestamp 1666464484
transform 1 0 30109 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_113
timestamp 1666464484
transform 1 0 37616 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_114
timestamp 1666464484
transform 1 0 41789 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_115
timestamp 1666464484
transform 1 0 41789 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_116
timestamp 1666464484
transform 1 0 50096 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_117
timestamp 1666464484
transform 1 0 50096 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_118
timestamp 1666464484
transform 1 0 41360 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_119
timestamp 1666464484
transform 1 0 41360 0 1 -1249
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_120
timestamp 1666464484
transform 1 0 40621 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_121
timestamp 1666464484
transform 1 0 40621 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_122
timestamp 1666464484
transform 1 0 48848 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_123
timestamp 1666464484
transform 1 0 48848 0 1 -1493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_124
timestamp 1666464484
transform 1 0 47600 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_125
timestamp 1666464484
transform 1 0 47600 0 1 -1737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_126
timestamp 1666464484
transform 1 0 46352 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_127
timestamp 1666464484
transform 1 0 46352 0 1 -1981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_128
timestamp 1666464484
transform 1 0 45104 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_129
timestamp 1666464484
transform 1 0 45104 0 1 -2225
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_130
timestamp 1666464484
transform 1 0 43856 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_131
timestamp 1666464484
transform 1 0 43856 0 1 -2469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_132
timestamp 1666464484
transform 1 0 44125 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_133
timestamp 1666464484
transform 1 0 44125 0 1 -2713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_134
timestamp 1666464484
transform 1 0 52592 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_135
timestamp 1666464484
transform 1 0 52592 0 1 -2713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_136
timestamp 1666464484
transform 1 0 43571 0 1 272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_137
timestamp 1666464484
transform 1 0 43571 0 1 -2713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_138
timestamp 1666464484
transform 1 0 42957 0 1 -3958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_139
timestamp 1666464484
transform 1 0 42957 0 1 -2957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_140
timestamp 1666464484
transform 1 0 51344 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_141
timestamp 1666464484
transform 1 0 51344 0 1 -2957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_142
timestamp 1666464484
transform 1 0 42608 0 1 1392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_143
timestamp 1666464484
transform 1 0 42608 0 1 -2957
box 0 0 1 1
<< properties >>
string FIXED_BBOX 3208 -3962 52705 1462
string GDS_END 7323320
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 7291268
<< end >>
