magic
tech sky130B
magscale 1 2
timestamp 1672550940
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 154114 700340 154120 700392
rect 154172 700380 154178 700392
rect 199378 700380 199384 700392
rect 154172 700352 199384 700380
rect 154172 700340 154178 700352
rect 199378 700340 199384 700352
rect 199436 700340 199442 700392
rect 202782 700340 202788 700392
rect 202840 700380 202846 700392
rect 203518 700380 203524 700392
rect 202840 700352 203524 700380
rect 202840 700340 202846 700352
rect 203518 700340 203524 700352
rect 203576 700340 203582 700392
rect 371878 700340 371884 700392
rect 371936 700380 371942 700392
rect 478506 700380 478512 700392
rect 371936 700352 478512 700380
rect 371936 700340 371942 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 206278 700312 206284 700324
rect 89220 700284 206284 700312
rect 89220 700272 89226 700284
rect 206278 700272 206284 700284
rect 206336 700272 206342 700324
rect 212534 700272 212540 700324
rect 212592 700312 212598 700324
rect 413646 700312 413652 700324
rect 212592 700284 413652 700312
rect 212592 700272 212598 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 418798 700272 418804 700324
rect 418856 700312 418862 700324
rect 429838 700312 429844 700324
rect 418856 700284 429844 700312
rect 418856 700272 418862 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 479518 700272 479524 700324
rect 479576 700312 479582 700324
rect 527174 700312 527180 700324
rect 479576 700284 527180 700312
rect 479576 700272 479582 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 8110 699660 8116 699712
rect 8168 699700 8174 699712
rect 10318 699700 10324 699712
rect 8168 699672 10324 699700
rect 8168 699660 8174 699672
rect 10318 699660 10324 699672
rect 10376 699660 10382 699712
rect 345658 699660 345664 699712
rect 345716 699700 345722 699712
rect 348786 699700 348792 699712
rect 345716 699672 348792 699700
rect 345716 699660 345722 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 558178 699660 558184 699712
rect 558236 699700 558242 699712
rect 559650 699700 559656 699712
rect 558236 699672 559656 699700
rect 558236 699660 558242 699672
rect 559650 699660 559656 699672
rect 559708 699660 559714 699712
rect 215294 697552 215300 697604
rect 215352 697592 215358 697604
rect 218974 697592 218980 697604
rect 215352 697564 218980 697592
rect 215352 697552 215358 697564
rect 218974 697552 218980 697564
rect 219032 697552 219038 697604
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 271138 696940 271144 696992
rect 271196 696980 271202 696992
rect 580166 696980 580172 696992
rect 271196 696952 580172 696980
rect 271196 696940 271202 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 23474 692044 23480 692096
rect 23532 692084 23538 692096
rect 219434 692084 219440 692096
rect 23532 692056 219440 692084
rect 23532 692044 23538 692056
rect 219434 692044 219440 692056
rect 219492 692044 219498 692096
rect 71774 690616 71780 690668
rect 71832 690656 71838 690668
rect 218054 690656 218060 690668
rect 71832 690628 218060 690656
rect 71832 690616 71838 690628
rect 218054 690616 218060 690628
rect 218112 690616 218118 690668
rect 136634 689256 136640 689308
rect 136692 689296 136698 689308
rect 216674 689296 216680 689308
rect 136692 689268 216680 689296
rect 136692 689256 136698 689268
rect 216674 689256 216680 689268
rect 216732 689256 216738 689308
rect 40034 687896 40040 687948
rect 40092 687936 40098 687948
rect 218146 687936 218152 687948
rect 40092 687908 218152 687936
rect 40092 687896 40098 687908
rect 218146 687896 218152 687908
rect 218204 687896 218210 687948
rect 104894 686468 104900 686520
rect 104952 686508 104958 686520
rect 216766 686508 216772 686520
rect 104952 686480 216772 686508
rect 104952 686468 104958 686480
rect 216766 686468 216772 686480
rect 216824 686468 216830 686520
rect 169754 685108 169760 685160
rect 169812 685148 169818 685160
rect 216858 685148 216864 685160
rect 169812 685120 216864 685148
rect 169812 685108 169818 685120
rect 216858 685108 216864 685120
rect 216916 685108 216922 685160
rect 166442 684904 166448 684956
rect 166500 684944 166506 684956
rect 249794 684944 249800 684956
rect 166500 684916 249800 684944
rect 166500 684904 166506 684916
rect 249794 684904 249800 684916
rect 249852 684904 249858 684956
rect 163958 684836 163964 684888
rect 164016 684876 164022 684888
rect 248414 684876 248420 684888
rect 164016 684848 248420 684876
rect 164016 684836 164022 684848
rect 248414 684836 248420 684848
rect 248472 684836 248478 684888
rect 159266 684768 159272 684820
rect 159324 684808 159330 684820
rect 244274 684808 244280 684820
rect 159324 684780 244280 684808
rect 159324 684768 159330 684780
rect 244274 684768 244280 684780
rect 244332 684768 244338 684820
rect 156874 684700 156880 684752
rect 156932 684740 156938 684752
rect 242894 684740 242900 684752
rect 156932 684712 242900 684740
rect 156932 684700 156938 684712
rect 242894 684700 242900 684712
rect 242952 684700 242958 684752
rect 154298 684632 154304 684684
rect 154356 684672 154362 684684
rect 240134 684672 240140 684684
rect 154356 684644 240140 684672
rect 154356 684632 154362 684644
rect 240134 684632 240140 684644
rect 240192 684632 240198 684684
rect 132954 684564 132960 684616
rect 133012 684604 133018 684616
rect 252554 684604 252560 684616
rect 133012 684576 252560 684604
rect 133012 684564 133018 684576
rect 252554 684564 252560 684576
rect 252612 684564 252618 684616
rect 118602 684496 118608 684548
rect 118660 684536 118666 684548
rect 241514 684536 241520 684548
rect 118660 684508 241520 684536
rect 118660 684496 118666 684508
rect 241514 684496 241520 684508
rect 241572 684496 241578 684548
rect 161382 684020 161388 684072
rect 161440 684060 161446 684072
rect 245654 684060 245660 684072
rect 161440 684032 245660 684060
rect 161440 684020 161446 684032
rect 245654 684020 245660 684032
rect 245712 684020 245718 684072
rect 142154 683952 142160 684004
rect 142212 683992 142218 684004
rect 242986 683992 242992 684004
rect 142212 683964 242992 683992
rect 142212 683952 142218 683964
rect 242986 683952 242992 683964
rect 243044 683952 243050 684004
rect 133874 683884 133880 683936
rect 133932 683924 133938 683936
rect 248506 683924 248512 683936
rect 133932 683896 248512 683924
rect 133932 683884 133938 683896
rect 248506 683884 248512 683896
rect 248564 683884 248570 683936
rect 130378 683816 130384 683868
rect 130436 683856 130442 683868
rect 247034 683856 247040 683868
rect 130436 683828 247040 683856
rect 130436 683816 130442 683828
rect 247034 683816 247040 683828
rect 247092 683816 247098 683868
rect 124214 683748 124220 683800
rect 124272 683788 124278 683800
rect 243078 683788 243084 683800
rect 124272 683760 243084 683788
rect 124272 683748 124278 683760
rect 243078 683748 243084 683760
rect 243136 683748 243142 683800
rect 111058 683680 111064 683732
rect 111116 683720 111122 683732
rect 241606 683720 241612 683732
rect 111116 683692 241612 683720
rect 111116 683680 111122 683692
rect 241606 683680 241612 683692
rect 241664 683680 241670 683732
rect 104250 683612 104256 683664
rect 104308 683652 104314 683664
rect 244366 683652 244372 683664
rect 104308 683624 244372 683652
rect 104308 683612 104314 683624
rect 244366 683612 244372 683624
rect 244424 683612 244430 683664
rect 97074 683544 97080 683596
rect 97132 683584 97138 683596
rect 238754 683584 238760 683596
rect 97132 683556 238760 683584
rect 97132 683544 97138 683556
rect 238754 683544 238760 683556
rect 238812 683544 238818 683596
rect 94682 683476 94688 683528
rect 94740 683516 94746 683528
rect 237650 683516 237656 683528
rect 94740 683488 237656 683516
rect 94740 683476 94746 683488
rect 237650 683476 237656 683488
rect 237708 683476 237714 683528
rect 92290 683408 92296 683460
rect 92348 683448 92354 683460
rect 235994 683448 236000 683460
rect 92348 683420 236000 683448
rect 92348 683408 92354 683420
rect 235994 683408 236000 683420
rect 236052 683408 236058 683460
rect 70762 683340 70768 683392
rect 70820 683380 70826 683392
rect 252646 683380 252652 683392
rect 70820 683352 252652 683380
rect 70820 683340 70826 683352
rect 252646 683340 252652 683352
rect 252704 683340 252710 683392
rect 44174 683272 44180 683324
rect 44232 683312 44238 683324
rect 241698 683312 241704 683324
rect 44232 683284 241704 683312
rect 44232 683272 44238 683284
rect 241698 683272 241704 683284
rect 241756 683272 241762 683324
rect 32490 683204 32496 683256
rect 32548 683244 32554 683256
rect 238846 683244 238852 683256
rect 32548 683216 238852 683244
rect 32548 683204 32554 683216
rect 238846 683204 238852 683216
rect 238904 683204 238910 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 202138 683176 202144 683188
rect 3476 683148 202144 683176
rect 3476 683136 3482 683148
rect 202138 683136 202144 683148
rect 202196 683136 202202 683188
rect 224218 683136 224224 683188
rect 224276 683176 224282 683188
rect 580166 683176 580172 683188
rect 224276 683148 580172 683176
rect 224276 683136 224282 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 61194 682864 61200 682916
rect 61252 682904 61258 682916
rect 146938 682904 146944 682916
rect 61252 682876 146944 682904
rect 61252 682864 61258 682876
rect 146938 682864 146944 682876
rect 146996 682864 147002 682916
rect 42058 682796 42064 682848
rect 42116 682836 42122 682848
rect 142154 682836 142160 682848
rect 42116 682808 142160 682836
rect 42116 682796 42122 682808
rect 142154 682796 142160 682808
rect 142212 682796 142218 682848
rect 85114 682728 85120 682780
rect 85172 682768 85178 682780
rect 137278 682768 137284 682780
rect 85172 682740 137284 682768
rect 85172 682728 85178 682740
rect 137278 682728 137284 682740
rect 137336 682728 137342 682780
rect 99282 682660 99288 682712
rect 99340 682700 99346 682712
rect 111058 682700 111064 682712
rect 99340 682672 111064 682700
rect 99340 682660 99346 682672
rect 111058 682660 111064 682672
rect 111116 682660 111122 682712
rect 106642 682592 106648 682644
rect 106700 682632 106706 682644
rect 130378 682632 130384 682644
rect 106700 682604 130384 682632
rect 106700 682592 106706 682604
rect 130378 682592 130384 682604
rect 130436 682592 130442 682644
rect 171042 682592 171048 682644
rect 171100 682632 171106 682644
rect 252738 682632 252744 682644
rect 171100 682604 252744 682632
rect 171100 682592 171106 682604
rect 252738 682592 252744 682604
rect 252796 682592 252802 682644
rect 101858 682524 101864 682576
rect 101916 682564 101922 682576
rect 124214 682564 124220 682576
rect 101916 682536 124220 682564
rect 101916 682524 101922 682536
rect 124214 682524 124220 682536
rect 124272 682524 124278 682576
rect 149698 682524 149704 682576
rect 149756 682564 149762 682576
rect 198182 682564 198188 682576
rect 149756 682536 198188 682564
rect 149756 682524 149762 682536
rect 198182 682524 198188 682536
rect 198240 682524 198246 682576
rect 108942 682456 108948 682508
rect 109000 682496 109006 682508
rect 133874 682496 133880 682508
rect 109000 682468 133880 682496
rect 109000 682456 109006 682468
rect 133874 682456 133880 682468
rect 133932 682456 133938 682508
rect 144822 682456 144828 682508
rect 144880 682496 144886 682508
rect 198274 682496 198280 682508
rect 144880 682468 198280 682496
rect 144880 682456 144886 682468
rect 198274 682456 198280 682468
rect 198332 682456 198338 682508
rect 142522 682388 142528 682440
rect 142580 682428 142586 682440
rect 197998 682428 198004 682440
rect 142580 682400 198004 682428
rect 142580 682388 142586 682400
rect 197998 682388 198004 682400
rect 198056 682388 198062 682440
rect 130562 682320 130568 682372
rect 130620 682360 130626 682372
rect 198090 682360 198096 682372
rect 130620 682332 198096 682360
rect 130620 682320 130626 682332
rect 198090 682320 198096 682332
rect 198148 682320 198154 682372
rect 44082 682252 44088 682304
rect 44140 682292 44146 682304
rect 168374 682292 168380 682304
rect 44140 682264 168380 682292
rect 44140 682252 44146 682264
rect 168374 682252 168380 682264
rect 168432 682252 168438 682304
rect 185578 682252 185584 682304
rect 185636 682292 185642 682304
rect 260834 682292 260840 682304
rect 185636 682264 260840 682292
rect 185636 682252 185642 682264
rect 260834 682252 260840 682264
rect 260892 682252 260898 682304
rect 65978 682184 65984 682236
rect 66036 682224 66042 682236
rect 100754 682224 100760 682236
rect 66036 682196 100760 682224
rect 66036 682184 66042 682196
rect 100754 682184 100760 682196
rect 100812 682184 100818 682236
rect 183186 682184 183192 682236
rect 183244 682224 183250 682236
rect 259730 682224 259736 682236
rect 183244 682196 259736 682224
rect 183244 682184 183250 682196
rect 259730 682184 259736 682196
rect 259788 682184 259794 682236
rect 58802 682116 58808 682168
rect 58860 682156 58866 682168
rect 107562 682156 107568 682168
rect 58860 682128 107568 682156
rect 58860 682116 58866 682128
rect 107562 682116 107568 682128
rect 107620 682116 107626 682168
rect 140130 682116 140136 682168
rect 140188 682156 140194 682168
rect 173802 682156 173808 682168
rect 140188 682128 173808 682156
rect 140188 682116 140194 682128
rect 173802 682116 173808 682128
rect 173860 682116 173866 682168
rect 178402 682116 178408 682168
rect 178460 682156 178466 682168
rect 256694 682156 256700 682168
rect 178460 682128 256700 682156
rect 178460 682116 178466 682128
rect 256694 682116 256700 682128
rect 256752 682116 256758 682168
rect 79962 682048 79968 682100
rect 80020 682088 80026 682100
rect 144270 682088 144276 682100
rect 80020 682060 144276 682088
rect 80020 682048 80026 682060
rect 144270 682048 144276 682060
rect 144328 682048 144334 682100
rect 180610 682048 180616 682100
rect 180668 682088 180674 682100
rect 258350 682088 258356 682100
rect 180668 682060 258356 682088
rect 180668 682048 180674 682060
rect 258350 682048 258356 682060
rect 258408 682048 258414 682100
rect 63402 681980 63408 682032
rect 63460 682020 63466 682032
rect 169754 682020 169760 682032
rect 63460 681992 169760 682020
rect 63460 681980 63466 681992
rect 169754 681980 169760 681992
rect 169812 681980 169818 682032
rect 176010 681980 176016 682032
rect 176068 682020 176074 682032
rect 255314 682020 255320 682032
rect 176068 681992 255320 682020
rect 176068 681980 176074 681992
rect 255314 681980 255320 681992
rect 255372 681980 255378 682032
rect 147306 681912 147312 681964
rect 147364 681952 147370 681964
rect 259546 681952 259552 681964
rect 147364 681924 259552 681952
rect 147364 681912 147370 681924
rect 259546 681912 259552 681924
rect 259604 681912 259610 681964
rect 25314 681844 25320 681896
rect 25372 681884 25378 681896
rect 60734 681884 60740 681896
rect 25372 681856 60740 681884
rect 25372 681844 25378 681856
rect 60734 681844 60740 681856
rect 60792 681844 60798 681896
rect 73062 681844 73068 681896
rect 73120 681884 73126 681896
rect 85482 681884 85488 681896
rect 73120 681856 85488 681884
rect 73120 681844 73126 681856
rect 85482 681844 85488 681856
rect 85540 681844 85546 681896
rect 128170 681844 128176 681896
rect 128228 681884 128234 681896
rect 249886 681884 249892 681896
rect 128228 681856 249892 681884
rect 128228 681844 128234 681856
rect 249886 681844 249892 681856
rect 249944 681844 249950 681896
rect 27522 681776 27528 681828
rect 27580 681816 27586 681828
rect 79042 681816 79048 681828
rect 27580 681788 79048 681816
rect 27580 681776 27586 681788
rect 79042 681776 79048 681788
rect 79100 681776 79106 681828
rect 125410 681776 125416 681828
rect 125468 681816 125474 681828
rect 247218 681816 247224 681828
rect 125468 681788 247224 681816
rect 125468 681776 125474 681788
rect 247218 681776 247224 681788
rect 247276 681776 247282 681828
rect 37182 681708 37188 681760
rect 37240 681748 37246 681760
rect 44174 681748 44180 681760
rect 37240 681720 44180 681748
rect 37240 681708 37246 681720
rect 44174 681708 44180 681720
rect 44232 681708 44238 681760
rect 87506 681708 87512 681760
rect 87564 681748 87570 681760
rect 98638 681748 98644 681760
rect 87564 681720 98644 681748
rect 87564 681708 87570 681720
rect 98638 681708 98644 681720
rect 98696 681708 98702 681760
rect 173618 681708 173624 681760
rect 173676 681748 173682 681760
rect 198366 681748 198372 681760
rect 173676 681720 198372 681748
rect 173676 681708 173682 681720
rect 198366 681708 198372 681720
rect 198424 681708 198430 681760
rect 168374 681300 168380 681352
rect 168432 681340 168438 681352
rect 243170 681340 243176 681352
rect 168432 681312 243176 681340
rect 168432 681300 168438 681312
rect 243170 681300 243176 681312
rect 243228 681300 243234 681352
rect 173802 681232 173808 681284
rect 173860 681272 173866 681284
rect 256786 681272 256792 681284
rect 173860 681244 256792 681272
rect 173860 681232 173866 681244
rect 256786 681232 256792 681244
rect 256844 681232 256850 681284
rect 146938 681164 146944 681216
rect 146996 681204 147002 681216
rect 249978 681204 249984 681216
rect 146996 681176 249984 681204
rect 146996 681164 147002 681176
rect 249978 681164 249984 681176
rect 250036 681164 250042 681216
rect 107562 681096 107568 681148
rect 107620 681136 107626 681148
rect 248690 681136 248696 681148
rect 107620 681108 248696 681136
rect 107620 681096 107626 681108
rect 248690 681096 248696 681108
rect 248748 681096 248754 681148
rect 100754 681028 100760 681080
rect 100812 681068 100818 681080
rect 251174 681068 251180 681080
rect 100812 681040 251180 681068
rect 100812 681028 100818 681040
rect 251174 681028 251180 681040
rect 251232 681028 251238 681080
rect 85482 680960 85488 681012
rect 85540 681000 85546 681012
rect 254210 681000 254216 681012
rect 85540 680972 254216 681000
rect 85540 680960 85546 680972
rect 254210 680960 254216 680972
rect 254268 680960 254274 681012
rect 123386 680824 123392 680876
rect 123444 680864 123450 680876
rect 245838 680864 245844 680876
rect 123444 680836 245844 680864
rect 123444 680824 123450 680836
rect 245838 680824 245844 680836
rect 245896 680824 245902 680876
rect 111426 680756 111432 680808
rect 111484 680796 111490 680808
rect 236178 680796 236184 680808
rect 111484 680768 236184 680796
rect 111484 680756 111490 680768
rect 236178 680756 236184 680768
rect 236236 680756 236242 680808
rect 82722 680688 82728 680740
rect 82780 680728 82786 680740
rect 256878 680728 256884 680740
rect 82780 680700 256884 680728
rect 82780 680688 82786 680700
rect 256878 680688 256884 680700
rect 256936 680688 256942 680740
rect 77938 680620 77944 680672
rect 77996 680660 78002 680672
rect 255406 680660 255412 680672
rect 77996 680632 255412 680660
rect 77996 680620 78002 680632
rect 255406 680620 255412 680632
rect 255464 680620 255470 680672
rect 68370 680552 68376 680604
rect 68428 680592 68434 680604
rect 252830 680592 252836 680604
rect 68428 680564 252836 680592
rect 68428 680552 68434 680564
rect 252830 680552 252836 680564
rect 252888 680552 252894 680604
rect 56410 680484 56416 680536
rect 56468 680524 56474 680536
rect 248598 680524 248604 680536
rect 56468 680496 248604 680524
rect 56468 680484 56474 680496
rect 248598 680484 248604 680496
rect 248656 680484 248662 680536
rect 49234 680416 49240 680468
rect 49292 680456 49298 680468
rect 245746 680456 245752 680468
rect 49292 680428 245752 680456
rect 49292 680416 49298 680428
rect 245746 680416 245752 680428
rect 245804 680416 245810 680468
rect 39666 680348 39672 680400
rect 39724 680388 39730 680400
rect 241790 680388 241796 680400
rect 39724 680360 241796 680388
rect 39724 680348 39730 680360
rect 241790 680348 241796 680360
rect 241848 680348 241854 680400
rect 137278 679668 137284 679720
rect 137336 679708 137342 679720
rect 258166 679708 258172 679720
rect 137336 679680 258172 679708
rect 137336 679668 137342 679680
rect 258166 679668 258172 679680
rect 258224 679668 258230 679720
rect 98638 679600 98644 679652
rect 98696 679640 98702 679652
rect 258258 679640 258264 679652
rect 98696 679612 258264 679640
rect 98696 679600 98702 679612
rect 258258 679600 258264 679612
rect 258316 679600 258322 679652
rect 89714 679396 89720 679448
rect 89772 679436 89778 679448
rect 89772 679408 93854 679436
rect 89772 679396 89778 679408
rect 93826 679028 93854 679408
rect 113818 679396 113824 679448
rect 113876 679396 113882 679448
rect 116026 679396 116032 679448
rect 116084 679396 116090 679448
rect 120994 679396 121000 679448
rect 121052 679436 121058 679448
rect 121052 679408 122834 679436
rect 121052 679396 121058 679408
rect 113836 679096 113864 679396
rect 116044 679164 116072 679396
rect 122806 679232 122834 679408
rect 135162 679396 135168 679448
rect 135220 679436 135226 679448
rect 135220 679408 142154 679436
rect 135220 679396 135226 679408
rect 142126 679300 142154 679408
rect 151906 679396 151912 679448
rect 151964 679436 151970 679448
rect 151964 679408 161474 679436
rect 151964 679396 151970 679408
rect 161446 679368 161474 679408
rect 187786 679396 187792 679448
rect 187844 679436 187850 679448
rect 234706 679436 234712 679448
rect 187844 679408 234712 679436
rect 187844 679396 187850 679408
rect 234706 679396 234712 679408
rect 234764 679396 234770 679448
rect 238938 679368 238944 679380
rect 161446 679340 238944 679368
rect 238938 679328 238944 679340
rect 238996 679328 239002 679380
rect 254026 679300 254032 679312
rect 142126 679272 254032 679300
rect 254026 679260 254032 679272
rect 254084 679260 254090 679312
rect 244550 679232 244556 679244
rect 122806 679204 244556 679232
rect 244550 679192 244556 679204
rect 244608 679192 244614 679244
rect 240318 679164 240324 679176
rect 116044 679136 240324 679164
rect 240318 679124 240324 679136
rect 240376 679124 240382 679176
rect 239030 679096 239036 679108
rect 113836 679068 239036 679096
rect 239030 679056 239036 679068
rect 239088 679056 239094 679108
rect 259638 679028 259644 679040
rect 93826 679000 259644 679028
rect 259638 678988 259644 679000
rect 259696 678988 259702 679040
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 20898 670732 20904 670744
rect 3568 670704 20904 670732
rect 3568 670692 3574 670704
rect 20898 670692 20904 670704
rect 20956 670692 20962 670744
rect 231118 670692 231124 670744
rect 231176 670732 231182 670744
rect 580166 670732 580172 670744
rect 231176 670704 580172 670732
rect 231176 670692 231182 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 11698 656928 11704 656940
rect 3476 656900 11704 656928
rect 3476 656888 3482 656900
rect 11698 656888 11704 656900
rect 11756 656888 11762 656940
rect 233878 643084 233884 643136
rect 233936 643124 233942 643136
rect 580166 643124 580172 643136
rect 233936 643096 580172 643124
rect 233936 643084 233942 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 208394 630640 208400 630692
rect 208452 630680 208458 630692
rect 580166 630680 580172 630692
rect 208452 630652 580172 630680
rect 208452 630640 208458 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 19978 618304 19984 618316
rect 3200 618276 19984 618304
rect 3200 618264 3206 618276
rect 19978 618264 19984 618276
rect 20036 618264 20042 618316
rect 222838 616836 222844 616888
rect 222896 616876 222902 616888
rect 580166 616876 580172 616888
rect 222896 616848 580172 616876
rect 222896 616836 222902 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 14458 605860 14464 605872
rect 3292 605832 14464 605860
rect 3292 605820 3298 605832
rect 14458 605820 14464 605832
rect 14516 605820 14522 605872
rect 228358 590656 228364 590708
rect 228416 590696 228422 590708
rect 579798 590696 579804 590708
rect 228416 590668 579804 590696
rect 228416 590656 228422 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 209774 588548 209780 588600
rect 209832 588588 209838 588600
rect 542354 588588 542360 588600
rect 209832 588560 542360 588588
rect 209832 588548 209838 588560
rect 542354 588548 542360 588560
rect 542412 588548 542418 588600
rect 211154 587120 211160 587172
rect 211212 587160 211218 587172
rect 462314 587160 462320 587172
rect 211212 587132 462320 587160
rect 211212 587120 211218 587132
rect 462314 587120 462320 587132
rect 462372 587120 462378 587172
rect 209866 585760 209872 585812
rect 209924 585800 209930 585812
rect 479518 585800 479524 585812
rect 209924 585772 479524 585800
rect 209924 585760 209930 585772
rect 479518 585760 479524 585772
rect 479576 585760 479582 585812
rect 551002 585148 551008 585200
rect 551060 585188 551066 585200
rect 557534 585188 557540 585200
rect 551060 585160 557540 585188
rect 551060 585148 551066 585160
rect 557534 585148 557540 585160
rect 557592 585148 557598 585200
rect 211246 584400 211252 584452
rect 211304 584440 211310 584452
rect 494054 584440 494060 584452
rect 211304 584412 494060 584440
rect 211304 584400 211310 584412
rect 494054 584400 494060 584412
rect 494112 584400 494118 584452
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 18598 579680 18604 579692
rect 3384 579652 18604 579680
rect 3384 579640 3390 579652
rect 18598 579640 18604 579652
rect 18656 579640 18662 579692
rect 562318 563048 562324 563100
rect 562376 563088 562382 563100
rect 580166 563088 580172 563100
rect 562376 563060 580172 563088
rect 562376 563048 562382 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 15838 553432 15844 553444
rect 3384 553404 15844 553432
rect 3384 553392 3390 553404
rect 15838 553392 15844 553404
rect 15896 553392 15902 553444
rect 406286 536800 406292 536852
rect 406344 536840 406350 536852
rect 416774 536840 416780 536852
rect 406344 536812 416780 536840
rect 406344 536800 406350 536812
rect 416774 536800 416780 536812
rect 416832 536800 416838 536852
rect 563698 536800 563704 536852
rect 563756 536840 563762 536852
rect 579890 536840 579896 536852
rect 563756 536812 579896 536840
rect 563756 536800 563762 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 270494 535440 270500 535492
rect 270552 535480 270558 535492
rect 416774 535480 416780 535492
rect 270552 535452 416780 535480
rect 270552 535440 270558 535452
rect 416774 535440 416780 535452
rect 416832 535440 416838 535492
rect 416038 532788 416044 532840
rect 416096 532828 416102 532840
rect 418062 532828 418068 532840
rect 416096 532800 418068 532828
rect 416096 532788 416102 532800
rect 418062 532788 418068 532800
rect 418120 532788 418126 532840
rect 280798 532720 280804 532772
rect 280856 532760 280862 532772
rect 417050 532760 417056 532772
rect 280856 532732 417056 532760
rect 280856 532720 280862 532732
rect 417050 532720 417056 532732
rect 417108 532720 417114 532772
rect 414658 530000 414664 530052
rect 414716 530040 414722 530052
rect 417418 530040 417424 530052
rect 414716 530012 417424 530040
rect 414716 530000 414722 530012
rect 417418 530000 417424 530012
rect 417476 530000 417482 530052
rect 279418 529932 279424 529984
rect 279476 529972 279482 529984
rect 417694 529972 417700 529984
rect 279476 529944 417700 529972
rect 279476 529932 279482 529944
rect 417694 529932 417700 529944
rect 417752 529932 417758 529984
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 7558 527184 7564 527196
rect 3016 527156 7564 527184
rect 3016 527144 3022 527156
rect 7558 527144 7564 527156
rect 7616 527144 7622 527196
rect 295978 527144 295984 527196
rect 296036 527184 296042 527196
rect 417694 527184 417700 527196
rect 296036 527156 417700 527184
rect 296036 527144 296042 527156
rect 417694 527144 417700 527156
rect 417752 527144 417758 527196
rect 565078 524424 565084 524476
rect 565136 524464 565142 524476
rect 580166 524464 580172 524476
rect 565136 524436 580172 524464
rect 565136 524424 565142 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 558270 510620 558276 510672
rect 558328 510660 558334 510672
rect 580166 510660 580172 510672
rect 558328 510632 580172 510660
rect 558328 510620 558334 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 277578 509260 277584 509312
rect 277636 509300 277642 509312
rect 417602 509300 417608 509312
rect 277636 509272 417608 509300
rect 277636 509260 277642 509272
rect 417602 509260 417608 509272
rect 417660 509260 417666 509312
rect 298738 507832 298744 507884
rect 298796 507872 298802 507884
rect 416774 507872 416780 507884
rect 298796 507844 416780 507872
rect 298796 507832 298802 507844
rect 416774 507832 416780 507844
rect 416832 507832 416838 507884
rect 213914 507084 213920 507136
rect 213972 507124 213978 507136
rect 345658 507124 345664 507136
rect 213972 507096 345664 507124
rect 213972 507084 213978 507096
rect 345658 507084 345664 507096
rect 345716 507084 345722 507136
rect 211338 505724 211344 505776
rect 211396 505764 211402 505776
rect 371878 505764 371884 505776
rect 211396 505736 371884 505764
rect 211396 505724 211402 505736
rect 371878 505724 371884 505736
rect 371936 505724 371942 505776
rect 214006 504364 214012 504416
rect 214064 504404 214070 504416
rect 331214 504404 331220 504416
rect 214064 504376 331220 504404
rect 214064 504364 214070 504376
rect 331214 504364 331220 504376
rect 331272 504364 331278 504416
rect 212626 502936 212632 502988
rect 212684 502976 212690 502988
rect 364334 502976 364340 502988
rect 212684 502948 364340 502976
rect 212684 502936 212690 502948
rect 364334 502936 364340 502948
rect 364392 502936 364398 502988
rect 212718 501576 212724 501628
rect 212776 501616 212782 501628
rect 396718 501616 396724 501628
rect 212776 501588 396724 501616
rect 212776 501576 212782 501588
rect 396718 501576 396724 501588
rect 396776 501576 396782 501628
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 20070 501004 20076 501016
rect 3384 500976 20076 501004
rect 3384 500964 3390 500976
rect 20070 500964 20076 500976
rect 20128 500964 20134 501016
rect 211430 500216 211436 500268
rect 211488 500256 211494 500268
rect 418798 500256 418804 500268
rect 211488 500228 418804 500256
rect 211488 500216 211494 500228
rect 418798 500216 418804 500228
rect 418856 500216 418862 500268
rect 205634 498788 205640 498840
rect 205692 498828 205698 498840
rect 558270 498828 558276 498840
rect 205692 498800 558276 498828
rect 205692 498788 205698 498800
rect 558270 498788 558276 498800
rect 558328 498788 558334 498840
rect 551922 498176 551928 498228
rect 551980 498216 551986 498228
rect 557534 498216 557540 498228
rect 551980 498188 557540 498216
rect 551980 498176 551986 498188
rect 557534 498176 557540 498188
rect 557592 498176 557598 498228
rect 476758 498040 476764 498092
rect 476816 498080 476822 498092
rect 480346 498080 480352 498092
rect 476816 498052 480352 498080
rect 476816 498040 476822 498052
rect 480346 498040 480352 498052
rect 480404 498040 480410 498092
rect 65242 497428 65248 497480
rect 65300 497468 65306 497480
rect 151078 497468 151084 497480
rect 65300 497440 151084 497468
rect 65300 497428 65306 497440
rect 151078 497428 151084 497440
rect 151136 497428 151142 497480
rect 276014 497224 276020 497276
rect 276072 497264 276078 497276
rect 485774 497264 485780 497276
rect 276072 497236 485780 497264
rect 276072 497224 276078 497236
rect 485774 497224 485780 497236
rect 485832 497224 485838 497276
rect 283558 497156 283564 497208
rect 283616 497196 283622 497208
rect 452654 497196 452660 497208
rect 283616 497168 452660 497196
rect 283616 497156 283622 497168
rect 452654 497156 452660 497168
rect 452712 497156 452718 497208
rect 262214 497088 262220 497140
rect 262272 497128 262278 497140
rect 436186 497128 436192 497140
rect 262272 497100 436192 497128
rect 262272 497088 262278 497100
rect 436186 497088 436192 497100
rect 436244 497088 436250 497140
rect 260926 497020 260932 497072
rect 260984 497060 260990 497072
rect 436094 497060 436100 497072
rect 260984 497032 436100 497060
rect 260984 497020 260990 497032
rect 436094 497020 436100 497032
rect 436152 497020 436158 497072
rect 457438 497020 457444 497072
rect 457496 497060 457502 497072
rect 473354 497060 473360 497072
rect 457496 497032 473360 497060
rect 457496 497020 457502 497032
rect 473354 497020 473360 497032
rect 473412 497020 473418 497072
rect 277486 496952 277492 497004
rect 277544 496992 277550 497004
rect 459554 496992 459560 497004
rect 277544 496964 459560 496992
rect 277544 496952 277550 496964
rect 459554 496952 459560 496964
rect 459612 496952 459618 497004
rect 464338 496952 464344 497004
rect 464396 496992 464402 497004
rect 476114 496992 476120 497004
rect 464396 496964 476120 496992
rect 464396 496952 464402 496964
rect 476114 496952 476120 496964
rect 476172 496952 476178 497004
rect 271874 496884 271880 496936
rect 271932 496924 271938 496936
rect 470778 496924 470784 496936
rect 271932 496896 470784 496924
rect 271932 496884 271938 496896
rect 470778 496884 470784 496896
rect 470836 496884 470842 496936
rect 475378 496884 475384 496936
rect 475436 496924 475442 496936
rect 483014 496924 483020 496936
rect 475436 496896 483020 496924
rect 475436 496884 475442 496896
rect 483014 496884 483020 496896
rect 483072 496884 483078 496936
rect 472618 496816 472624 496868
rect 472676 496856 472682 496868
rect 477494 496856 477500 496868
rect 472676 496828 477500 496856
rect 472676 496816 472682 496828
rect 477494 496816 477500 496828
rect 477552 496816 477558 496868
rect 269114 496136 269120 496188
rect 269172 496176 269178 496188
rect 448514 496176 448520 496188
rect 269172 496148 448520 496176
rect 269172 496136 269178 496148
rect 448514 496136 448520 496148
rect 448572 496136 448578 496188
rect 274634 496068 274640 496120
rect 274692 496108 274698 496120
rect 455414 496108 455420 496120
rect 274692 496080 455420 496108
rect 274692 496068 274698 496080
rect 455414 496068 455420 496080
rect 455472 496068 455478 496120
rect 262306 494708 262312 494760
rect 262364 494748 262370 494760
rect 437474 494748 437480 494760
rect 262364 494720 437480 494748
rect 262364 494708 262370 494720
rect 437474 494708 437480 494720
rect 437532 494708 437538 494760
rect 273254 493280 273260 493332
rect 273312 493320 273318 493332
rect 454034 493320 454040 493332
rect 273312 493292 454040 493320
rect 273312 493280 273318 493292
rect 454034 493280 454040 493292
rect 454092 493280 454098 493332
rect 215386 491988 215392 492040
rect 215444 492028 215450 492040
rect 282914 492028 282920 492040
rect 215444 492000 282920 492028
rect 215444 491988 215450 492000
rect 282914 491988 282920 492000
rect 282972 491988 282978 492040
rect 276106 491920 276112 491972
rect 276164 491960 276170 491972
rect 458266 491960 458272 491972
rect 276164 491932 458272 491960
rect 276164 491920 276170 491932
rect 458266 491920 458272 491932
rect 458324 491920 458330 491972
rect 274726 490560 274732 490612
rect 274784 490600 274790 490612
rect 456886 490600 456892 490612
rect 274784 490572 456892 490600
rect 274784 490560 274790 490572
rect 456886 490560 456892 490572
rect 456944 490560 456950 490612
rect 276198 489200 276204 489252
rect 276256 489240 276262 489252
rect 456794 489240 456800 489252
rect 276256 489212 456800 489240
rect 276256 489200 276262 489212
rect 456794 489200 456800 489212
rect 456852 489200 456858 489252
rect 205726 489132 205732 489184
rect 205784 489172 205790 489184
rect 562318 489172 562324 489184
rect 205784 489144 562324 489172
rect 205784 489132 205790 489144
rect 562318 489132 562324 489144
rect 562376 489132 562382 489184
rect 262398 487772 262404 487824
rect 262456 487812 262462 487824
rect 443086 487812 443092 487824
rect 262456 487784 443092 487812
rect 262456 487772 262462 487784
rect 443086 487772 443092 487784
rect 443144 487772 443150 487824
rect 266446 486412 266452 486464
rect 266504 486452 266510 486464
rect 441614 486452 441620 486464
rect 266504 486424 441620 486452
rect 266504 486412 266510 486424
rect 441614 486412 441620 486424
rect 441672 486412 441678 486464
rect 226978 484372 226984 484424
rect 227036 484412 227042 484424
rect 580166 484412 580172 484424
rect 227036 484384 580172 484412
rect 227036 484372 227042 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 263594 483624 263600 483676
rect 263652 483664 263658 483676
rect 438854 483664 438860 483676
rect 263652 483636 438860 483664
rect 263652 483624 263658 483636
rect 438854 483624 438860 483636
rect 438912 483624 438918 483676
rect 209958 482332 209964 482384
rect 210016 482372 210022 482384
rect 224218 482372 224224 482384
rect 210016 482344 224224 482372
rect 210016 482332 210022 482344
rect 224218 482332 224224 482344
rect 224276 482332 224282 482384
rect 3510 482264 3516 482316
rect 3568 482304 3574 482316
rect 223574 482304 223580 482316
rect 3568 482276 223580 482304
rect 3568 482264 3574 482276
rect 223574 482264 223580 482276
rect 223632 482264 223638 482316
rect 271966 482264 271972 482316
rect 272024 482304 272030 482316
rect 467834 482304 467840 482316
rect 272024 482276 467840 482304
rect 272024 482264 272030 482276
rect 467834 482264 467840 482276
rect 467892 482264 467898 482316
rect 3418 480972 3424 481024
rect 3476 481012 3482 481024
rect 222194 481012 222200 481024
rect 3476 480984 222200 481012
rect 3476 480972 3482 480984
rect 222194 480972 222200 480984
rect 222252 480972 222258 481024
rect 270586 480972 270592 481024
rect 270644 481012 270650 481024
rect 465074 481012 465080 481024
rect 270644 480984 465080 481012
rect 270644 480972 270650 480984
rect 465074 480972 465080 480984
rect 465132 480972 465138 481024
rect 207014 480904 207020 480956
rect 207072 480944 207078 480956
rect 580258 480944 580264 480956
rect 207072 480916 580264 480944
rect 207072 480904 207078 480916
rect 580258 480904 580264 480916
rect 580316 480904 580322 480956
rect 19978 479544 19984 479596
rect 20036 479584 20042 479596
rect 220814 479584 220820 479596
rect 20036 479556 220820 479584
rect 20036 479544 20042 479556
rect 220814 479544 220820 479556
rect 220872 479544 220878 479596
rect 269206 479544 269212 479596
rect 269264 479584 269270 479596
rect 460934 479584 460940 479596
rect 269264 479556 460940 479584
rect 269264 479544 269270 479556
rect 460934 479544 460940 479556
rect 460992 479544 460998 479596
rect 205818 479476 205824 479528
rect 205876 479516 205882 479528
rect 565078 479516 565084 479528
rect 205876 479488 565084 479516
rect 205876 479476 205882 479488
rect 565078 479476 565084 479488
rect 565136 479476 565142 479528
rect 208486 478184 208492 478236
rect 208544 478224 208550 478236
rect 271138 478224 271144 478236
rect 208544 478196 271144 478224
rect 208544 478184 208550 478196
rect 271138 478184 271144 478196
rect 271196 478184 271202 478236
rect 21358 478116 21364 478168
rect 21416 478156 21422 478168
rect 220906 478156 220912 478168
rect 21416 478128 220912 478156
rect 21416 478116 21422 478128
rect 220906 478116 220912 478128
rect 220964 478116 220970 478168
rect 269298 478116 269304 478168
rect 269356 478156 269362 478168
rect 462314 478156 462320 478168
rect 269356 478128 462320 478156
rect 269356 478116 269362 478128
rect 462314 478116 462320 478128
rect 462372 478116 462378 478168
rect 206278 476892 206284 476944
rect 206336 476932 206342 476944
rect 218238 476932 218244 476944
rect 206336 476904 218244 476932
rect 206336 476892 206342 476904
rect 218238 476892 218244 476904
rect 218296 476892 218302 476944
rect 214098 476824 214104 476876
rect 214156 476864 214162 476876
rect 266354 476864 266360 476876
rect 214156 476836 266360 476864
rect 214156 476824 214162 476836
rect 266354 476824 266360 476836
rect 266412 476824 266418 476876
rect 22094 476756 22100 476808
rect 22152 476796 22158 476808
rect 236270 476796 236276 476808
rect 22152 476768 236276 476796
rect 22152 476756 22158 476768
rect 236270 476756 236276 476768
rect 236328 476756 236334 476808
rect 267734 476756 267740 476808
rect 267792 476796 267798 476808
rect 458174 476796 458180 476808
rect 267792 476768 458180 476796
rect 267792 476756 267798 476768
rect 458174 476756 458180 476768
rect 458232 476756 458238 476808
rect 266354 475328 266360 475380
rect 266412 475368 266418 475380
rect 454678 475368 454684 475380
rect 266412 475340 454684 475368
rect 266412 475328 266418 475340
rect 454678 475328 454684 475340
rect 454736 475328 454742 475380
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 223666 474756 223672 474768
rect 3476 474728 223672 474756
rect 3476 474716 3482 474728
rect 223666 474716 223672 474728
rect 223724 474716 223730 474768
rect 20070 474036 20076 474088
rect 20128 474076 20134 474088
rect 223758 474076 223764 474088
rect 20128 474048 223764 474076
rect 20128 474036 20134 474048
rect 223758 474036 223764 474048
rect 223816 474036 223822 474088
rect 264974 474036 264980 474088
rect 265032 474076 265038 474088
rect 452746 474076 452752 474088
rect 265032 474048 452752 474076
rect 265032 474036 265038 474048
rect 452746 474036 452752 474048
rect 452804 474036 452810 474088
rect 205910 473968 205916 474020
rect 205968 474008 205974 474020
rect 563698 474008 563704 474020
rect 205968 473980 563704 474008
rect 205968 473968 205974 473980
rect 563698 473968 563704 473980
rect 563756 473968 563762 474020
rect 214190 472676 214196 472728
rect 214248 472716 214254 472728
rect 299474 472716 299480 472728
rect 214248 472688 299480 472716
rect 214248 472676 214254 472688
rect 299474 472676 299480 472688
rect 299532 472676 299538 472728
rect 15838 472608 15844 472660
rect 15896 472648 15902 472660
rect 222286 472648 222292 472660
rect 15896 472620 222292 472648
rect 15896 472608 15902 472620
rect 222286 472608 222292 472620
rect 222344 472608 222350 472660
rect 263686 472608 263692 472660
rect 263744 472648 263750 472660
rect 449986 472648 449992 472660
rect 263744 472620 449992 472648
rect 263744 472608 263750 472620
rect 449986 472608 449992 472620
rect 450044 472608 450050 472660
rect 14458 471248 14464 471300
rect 14516 471288 14522 471300
rect 220998 471288 221004 471300
rect 14516 471260 221004 471288
rect 14516 471248 14522 471260
rect 220998 471248 221004 471260
rect 221056 471248 221062 471300
rect 270678 471248 270684 471300
rect 270736 471288 270742 471300
rect 451366 471288 451372 471300
rect 270736 471260 451372 471288
rect 270736 471248 270742 471260
rect 451366 471248 451372 471260
rect 451424 471248 451430 471300
rect 204254 470568 204260 470620
rect 204312 470608 204318 470620
rect 579982 470608 579988 470620
rect 204312 470580 579988 470608
rect 204312 470568 204318 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 207106 469888 207112 469940
rect 207164 469928 207170 469940
rect 228358 469928 228364 469940
rect 207164 469900 228364 469928
rect 207164 469888 207170 469900
rect 228358 469888 228364 469900
rect 228416 469888 228422 469940
rect 270770 469888 270776 469940
rect 270828 469928 270834 469940
rect 449894 469928 449900 469940
rect 270828 469900 449900 469928
rect 270828 469888 270834 469900
rect 449894 469888 449900 469900
rect 449952 469888 449958 469940
rect 11698 469820 11704 469872
rect 11756 469860 11762 469872
rect 219526 469860 219532 469872
rect 11756 469832 219532 469860
rect 11756 469820 11762 469832
rect 219526 469820 219532 469832
rect 219584 469820 219590 469872
rect 273346 469820 273352 469872
rect 273404 469860 273410 469872
rect 464338 469860 464344 469872
rect 273404 469832 464344 469860
rect 273404 469820 273410 469832
rect 464338 469820 464344 469832
rect 464396 469820 464402 469872
rect 204346 468528 204352 468580
rect 204404 468568 204410 468580
rect 226978 468568 226984 468580
rect 204404 468540 226984 468568
rect 204404 468528 204410 468540
rect 226978 468528 226984 468540
rect 227036 468528 227042 468580
rect 267826 468528 267832 468580
rect 267884 468568 267890 468580
rect 447226 468568 447232 468580
rect 267884 468540 447232 468568
rect 267884 468528 267890 468540
rect 447226 468528 447232 468540
rect 447284 468528 447290 468580
rect 10318 468460 10324 468512
rect 10376 468500 10382 468512
rect 219618 468500 219624 468512
rect 10376 468472 219624 468500
rect 10376 468460 10382 468472
rect 219618 468460 219624 468472
rect 219676 468460 219682 468512
rect 273438 468460 273444 468512
rect 273496 468500 273502 468512
rect 457438 468500 457444 468512
rect 273496 468472 457444 468500
rect 273496 468460 273502 468472
rect 457438 468460 457444 468472
rect 457496 468460 457502 468512
rect 208578 467168 208584 467220
rect 208636 467208 208642 467220
rect 233878 467208 233884 467220
rect 208636 467180 233884 467208
rect 208636 467168 208642 467180
rect 233878 467168 233884 467180
rect 233936 467168 233942 467220
rect 261018 467168 261024 467220
rect 261076 467208 261082 467220
rect 298738 467208 298744 467220
rect 261076 467180 298744 467208
rect 261076 467168 261082 467180
rect 298738 467168 298744 467180
rect 298796 467168 298802 467220
rect 7558 467100 7564 467152
rect 7616 467140 7622 467152
rect 222378 467140 222384 467152
rect 7616 467112 222384 467140
rect 7616 467100 7622 467112
rect 222378 467100 222384 467112
rect 222436 467100 222442 467152
rect 276290 467100 276296 467152
rect 276348 467140 276354 467152
rect 475378 467140 475384 467152
rect 276348 467112 475384 467140
rect 276348 467100 276354 467112
rect 475378 467100 475384 467112
rect 475436 467100 475442 467152
rect 198918 466828 198924 466880
rect 198976 466868 198982 466880
rect 577682 466868 577688 466880
rect 198976 466840 577688 466868
rect 198976 466828 198982 466840
rect 577682 466828 577688 466840
rect 577740 466828 577746 466880
rect 198826 466760 198832 466812
rect 198884 466800 198890 466812
rect 577866 466800 577872 466812
rect 198884 466772 577872 466800
rect 198884 466760 198890 466772
rect 577866 466760 577872 466772
rect 577924 466760 577930 466812
rect 198734 466692 198740 466744
rect 198792 466732 198798 466744
rect 577958 466732 577964 466744
rect 198792 466704 577964 466732
rect 198792 466692 198798 466704
rect 577958 466692 577964 466704
rect 578016 466692 578022 466744
rect 200114 466624 200120 466676
rect 200172 466664 200178 466676
rect 580534 466664 580540 466676
rect 200172 466636 580540 466664
rect 200172 466624 200178 466636
rect 580534 466624 580540 466636
rect 580592 466624 580598 466676
rect 197630 466556 197636 466608
rect 197688 466596 197694 466608
rect 577774 466596 577780 466608
rect 197688 466568 577780 466596
rect 197688 466556 197694 466568
rect 577774 466556 577780 466568
rect 577832 466556 577838 466608
rect 196066 466488 196072 466540
rect 196124 466528 196130 466540
rect 577498 466528 577504 466540
rect 196124 466500 577504 466528
rect 196124 466488 196130 466500
rect 577498 466488 577504 466500
rect 577556 466488 577562 466540
rect 196158 466420 196164 466472
rect 196216 466460 196222 466472
rect 580258 466460 580264 466472
rect 196216 466432 580264 466460
rect 196216 466420 196222 466432
rect 580258 466420 580264 466432
rect 580316 466420 580322 466472
rect 269390 465808 269396 465860
rect 269448 465848 269454 465860
rect 280798 465848 280804 465860
rect 269448 465820 280804 465848
rect 269448 465808 269454 465820
rect 280798 465808 280804 465820
rect 280856 465808 280862 465860
rect 18598 465740 18604 465792
rect 18656 465780 18662 465792
rect 222470 465780 222476 465792
rect 18656 465752 222476 465780
rect 18656 465740 18662 465752
rect 222470 465740 222476 465752
rect 222528 465740 222534 465792
rect 274818 465740 274824 465792
rect 274876 465780 274882 465792
rect 472618 465780 472624 465792
rect 274876 465752 472624 465780
rect 274876 465740 274882 465752
rect 472618 465740 472624 465752
rect 472676 465740 472682 465792
rect 210050 465672 210056 465724
rect 210108 465712 210114 465724
rect 558178 465712 558184 465724
rect 210108 465684 558184 465712
rect 210108 465672 210114 465684
rect 558178 465672 558184 465684
rect 558236 465672 558242 465724
rect 160738 465468 160744 465520
rect 160796 465508 160802 465520
rect 367094 465508 367100 465520
rect 160796 465480 367100 465508
rect 160796 465468 160802 465480
rect 367094 465468 367100 465480
rect 367152 465468 367158 465520
rect 161014 465400 161020 465452
rect 161072 465440 161078 465452
rect 370130 465440 370136 465452
rect 161072 465412 370136 465440
rect 161072 465400 161078 465412
rect 370130 465400 370136 465412
rect 370188 465400 370194 465452
rect 160922 465332 160928 465384
rect 160980 465372 160986 465384
rect 372614 465372 372620 465384
rect 160980 465344 372620 465372
rect 160980 465332 160986 465344
rect 372614 465332 372620 465344
rect 372672 465332 372678 465384
rect 160830 465264 160836 465316
rect 160888 465304 160894 465316
rect 375374 465304 375380 465316
rect 160888 465276 375380 465304
rect 160888 465264 160894 465276
rect 375374 465264 375380 465276
rect 375432 465264 375438 465316
rect 14642 465196 14648 465248
rect 14700 465236 14706 465248
rect 231946 465236 231952 465248
rect 14700 465208 231952 465236
rect 14700 465196 14706 465208
rect 231946 465196 231952 465208
rect 232004 465196 232010 465248
rect 197446 465128 197452 465180
rect 197504 465168 197510 465180
rect 577590 465168 577596 465180
rect 197504 465140 577596 465168
rect 197504 465128 197510 465140
rect 577590 465128 577596 465140
rect 577648 465128 577654 465180
rect 197538 465060 197544 465112
rect 197596 465100 197602 465112
rect 580350 465100 580356 465112
rect 197596 465072 580356 465100
rect 197596 465060 197602 465072
rect 580350 465060 580356 465072
rect 580408 465060 580414 465112
rect 169018 464584 169024 464636
rect 169076 464624 169082 464636
rect 327350 464624 327356 464636
rect 169076 464596 327356 464624
rect 169076 464584 169082 464596
rect 327350 464584 327356 464596
rect 327408 464584 327414 464636
rect 316310 464516 316316 464568
rect 316368 464556 316374 464568
rect 395338 464556 395344 464568
rect 316368 464528 395344 464556
rect 316368 464516 316374 464528
rect 395338 464516 395344 464528
rect 395396 464516 395402 464568
rect 199378 464448 199384 464500
rect 199436 464488 199442 464500
rect 216950 464488 216956 464500
rect 199436 464460 216956 464488
rect 199436 464448 199442 464460
rect 216950 464448 216956 464460
rect 217008 464448 217014 464500
rect 302234 464448 302240 464500
rect 302292 464488 302298 464500
rect 394050 464488 394056 464500
rect 302292 464460 394056 464488
rect 302292 464448 302298 464460
rect 394050 464448 394056 464460
rect 394108 464448 394114 464500
rect 208670 464380 208676 464432
rect 208728 464420 208734 464432
rect 231118 464420 231124 464432
rect 208728 464392 231124 464420
rect 208728 464380 208734 464392
rect 231118 464380 231124 464392
rect 231176 464380 231182 464432
rect 267918 464380 267924 464432
rect 267976 464420 267982 464432
rect 416038 464420 416044 464432
rect 267976 464392 416044 464420
rect 267976 464380 267982 464392
rect 416038 464380 416044 464392
rect 416096 464380 416102 464432
rect 4798 464312 4804 464364
rect 4856 464352 4862 464364
rect 221090 464352 221096 464364
rect 4856 464324 221096 464352
rect 4856 464312 4862 464324
rect 221090 464312 221096 464324
rect 221148 464312 221154 464364
rect 266538 464312 266544 464364
rect 266596 464352 266602 464364
rect 445754 464352 445760 464364
rect 266596 464324 445760 464352
rect 266596 464312 266602 464324
rect 445754 464312 445760 464324
rect 445812 464312 445818 464364
rect 320358 464244 320364 464296
rect 320416 464284 320422 464296
rect 406194 464284 406200 464296
rect 320416 464256 406200 464284
rect 320416 464244 320422 464256
rect 406194 464244 406200 464256
rect 406252 464244 406258 464296
rect 166718 464176 166724 464228
rect 166776 464216 166782 464228
rect 331490 464216 331496 464228
rect 166776 464188 331496 464216
rect 166776 464176 166782 464188
rect 331490 464176 331496 464188
rect 331548 464176 331554 464228
rect 166350 464108 166356 464160
rect 166408 464148 166414 464160
rect 333974 464148 333980 464160
rect 166408 464120 333980 464148
rect 166408 464108 166414 464120
rect 333974 464108 333980 464120
rect 334032 464108 334038 464160
rect 166810 464040 166816 464092
rect 166868 464080 166874 464092
rect 336734 464080 336740 464092
rect 166868 464052 336740 464080
rect 166868 464040 166874 464052
rect 336734 464040 336740 464052
rect 336792 464040 336798 464092
rect 166534 463972 166540 464024
rect 166592 464012 166598 464024
rect 341150 464012 341156 464024
rect 166592 463984 341156 464012
rect 166592 463972 166598 463984
rect 341150 463972 341156 463984
rect 341208 463972 341214 464024
rect 166442 463904 166448 463956
rect 166500 463944 166506 463956
rect 343634 463944 343640 463956
rect 166500 463916 343640 463944
rect 166500 463904 166506 463916
rect 343634 463904 343640 463916
rect 343692 463904 343698 463956
rect 166258 463836 166264 463888
rect 166316 463876 166322 463888
rect 346578 463876 346584 463888
rect 166316 463848 346584 463876
rect 166316 463836 166322 463848
rect 346578 463836 346584 463848
rect 346636 463836 346642 463888
rect 171778 463768 171784 463820
rect 171836 463808 171842 463820
rect 380894 463808 380900 463820
rect 171836 463780 380900 463808
rect 171836 463768 171842 463780
rect 380894 463768 380900 463780
rect 380952 463768 380958 463820
rect 199010 463700 199016 463752
rect 199068 463740 199074 463752
rect 580442 463740 580448 463752
rect 199068 463712 580448 463740
rect 199068 463700 199074 463712
rect 580442 463700 580448 463712
rect 580500 463700 580506 463752
rect 174630 463292 174636 463344
rect 174688 463332 174694 463344
rect 378134 463332 378140 463344
rect 174688 463304 378140 463332
rect 174688 463292 174694 463304
rect 378134 463292 378140 463304
rect 378192 463292 378198 463344
rect 202138 463224 202144 463276
rect 202196 463264 202202 463276
rect 219710 463264 219716 463276
rect 202196 463236 219716 463264
rect 202196 463224 202202 463236
rect 219710 463224 219716 463236
rect 219768 463224 219774 463276
rect 266630 463224 266636 463276
rect 266688 463264 266694 463276
rect 279418 463264 279424 463276
rect 266688 463236 279424 463264
rect 266688 463224 266694 463236
rect 279418 463224 279424 463236
rect 279476 463224 279482 463276
rect 159726 463156 159732 463208
rect 159784 463196 159790 463208
rect 294138 463196 294144 463208
rect 159784 463168 294144 463196
rect 159784 463156 159790 463168
rect 294138 463156 294144 463168
rect 294196 463156 294202 463208
rect 349246 463156 349252 463208
rect 349304 463196 349310 463208
rect 407850 463196 407856 463208
rect 349304 463168 407856 463196
rect 349304 463156 349310 463168
rect 407850 463156 407856 463168
rect 407908 463156 407914 463208
rect 159634 463088 159640 463140
rect 159692 463128 159698 463140
rect 298186 463128 298192 463140
rect 159692 463100 298192 463128
rect 159692 463088 159698 463100
rect 298186 463088 298192 463100
rect 298244 463088 298250 463140
rect 346486 463088 346492 463140
rect 346544 463128 346550 463140
rect 410610 463128 410616 463140
rect 346544 463100 410616 463128
rect 346544 463088 346550 463100
rect 410610 463088 410616 463100
rect 410668 463088 410674 463140
rect 159358 463020 159364 463072
rect 159416 463060 159422 463072
rect 302326 463060 302332 463072
rect 159416 463032 302332 463060
rect 159416 463020 159422 463032
rect 302326 463020 302332 463032
rect 302384 463020 302390 463072
rect 342254 463020 342260 463072
rect 342312 463060 342318 463072
rect 410702 463060 410708 463072
rect 342312 463032 410708 463060
rect 342312 463020 342318 463032
rect 410702 463020 410708 463032
rect 410760 463020 410766 463072
rect 167730 462952 167736 463004
rect 167788 462992 167794 463004
rect 233510 462992 233516 463004
rect 167788 462964 233516 462992
rect 167788 462952 167794 462964
rect 233510 462952 233516 462964
rect 233568 462952 233574 463004
rect 261110 462952 261116 463004
rect 261168 462992 261174 463004
rect 447134 462992 447140 463004
rect 261168 462964 447140 462992
rect 261168 462952 261174 462964
rect 447134 462952 447140 462964
rect 447192 462952 447198 463004
rect 159542 462884 159548 462936
rect 159600 462924 159606 462936
rect 306374 462924 306380 462936
rect 159600 462896 306380 462924
rect 159600 462884 159606 462896
rect 306374 462884 306380 462896
rect 306432 462884 306438 462936
rect 336826 462884 336832 462936
rect 336884 462924 336890 462936
rect 407758 462924 407764 462936
rect 336884 462896 407764 462924
rect 336884 462884 336890 462896
rect 407758 462884 407764 462896
rect 407816 462884 407822 462936
rect 309134 462816 309140 462868
rect 309192 462856 309198 462868
rect 395430 462856 395436 462868
rect 309192 462828 395436 462856
rect 309192 462816 309198 462828
rect 395430 462816 395436 462828
rect 395488 462816 395494 462868
rect 159450 462748 159456 462800
rect 159508 462788 159514 462800
rect 314654 462788 314660 462800
rect 159508 462760 314660 462788
rect 159508 462748 159514 462760
rect 314654 462748 314660 462760
rect 314712 462748 314718 462800
rect 330110 462748 330116 462800
rect 330168 462788 330174 462800
rect 408034 462788 408040 462800
rect 330168 462760 408040 462788
rect 330168 462748 330174 462760
rect 408034 462748 408040 462760
rect 408092 462748 408098 462800
rect 162118 462680 162124 462732
rect 162176 462720 162182 462732
rect 317414 462720 317420 462732
rect 162176 462692 317420 462720
rect 162176 462680 162182 462692
rect 317414 462680 317420 462692
rect 317472 462680 317478 462732
rect 323118 462680 323124 462732
rect 323176 462720 323182 462732
rect 404998 462720 405004 462732
rect 323176 462692 405004 462720
rect 323176 462680 323182 462692
rect 404998 462680 405004 462692
rect 405056 462680 405062 462732
rect 161106 462612 161112 462664
rect 161164 462652 161170 462664
rect 310514 462652 310520 462664
rect 161164 462624 310520 462652
rect 161164 462612 161170 462624
rect 310514 462612 310520 462624
rect 310572 462612 310578 462664
rect 339494 462612 339500 462664
rect 339552 462652 339558 462664
rect 407942 462652 407948 462664
rect 339552 462624 407948 462652
rect 339552 462612 339558 462624
rect 407942 462612 407948 462624
rect 408000 462612 408006 462664
rect 174538 462544 174544 462596
rect 174596 462584 174602 462596
rect 375466 462584 375472 462596
rect 174596 462556 375472 462584
rect 174596 462544 174602 462556
rect 375466 462544 375472 462556
rect 375524 462544 375530 462596
rect 163682 462476 163688 462528
rect 163740 462516 163746 462528
rect 351914 462516 351920 462528
rect 163740 462488 351920 462516
rect 163740 462476 163746 462488
rect 351914 462476 351920 462488
rect 351972 462476 351978 462528
rect 354766 462476 354772 462528
rect 354824 462516 354830 462528
rect 410794 462516 410800 462528
rect 354824 462488 410800 462516
rect 354824 462476 354830 462488
rect 410794 462476 410800 462488
rect 410852 462476 410858 462528
rect 14550 462408 14556 462460
rect 14608 462448 14614 462460
rect 232038 462448 232044 462460
rect 14608 462420 232044 462448
rect 14608 462408 14614 462420
rect 232038 462408 232044 462420
rect 232096 462408 232102 462460
rect 304994 462408 305000 462460
rect 305052 462448 305058 462460
rect 403618 462448 403624 462460
rect 305052 462420 403624 462448
rect 305052 462408 305058 462420
rect 403618 462408 403624 462420
rect 403676 462408 403682 462460
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 225138 462380 225144 462392
rect 3292 462352 225144 462380
rect 3292 462340 3298 462352
rect 225138 462340 225144 462352
rect 225196 462340 225202 462392
rect 298278 462340 298284 462392
rect 298336 462380 298342 462392
rect 416038 462380 416044 462392
rect 298336 462352 416044 462380
rect 298336 462340 298342 462352
rect 416038 462340 416044 462352
rect 416096 462340 416102 462392
rect 177298 461932 177304 461984
rect 177356 461972 177362 461984
rect 342346 461972 342352 461984
rect 177356 461944 342352 461972
rect 177356 461932 177362 461944
rect 342346 461932 342352 461944
rect 342404 461932 342410 461984
rect 167914 461864 167920 461916
rect 167972 461904 167978 461916
rect 229094 461904 229100 461916
rect 167972 461876 229100 461904
rect 167972 461864 167978 461876
rect 229094 461864 229100 461876
rect 229152 461864 229158 461916
rect 195974 461796 195980 461848
rect 196032 461836 196038 461848
rect 196158 461836 196164 461848
rect 196032 461808 196164 461836
rect 196032 461796 196038 461808
rect 196158 461796 196164 461808
rect 196216 461796 196222 461848
rect 203518 461796 203524 461848
rect 203576 461836 203582 461848
rect 215570 461836 215576 461848
rect 203576 461808 215576 461836
rect 203576 461796 203582 461808
rect 215570 461796 215576 461808
rect 215628 461796 215634 461848
rect 161198 461728 161204 461780
rect 161256 461768 161262 461780
rect 289998 461768 290004 461780
rect 161256 461740 290004 461768
rect 161256 461728 161262 461740
rect 289998 461728 290004 461740
rect 290056 461728 290062 461780
rect 313274 461728 313280 461780
rect 313332 461768 313338 461780
rect 395522 461768 395528 461780
rect 313332 461740 395528 461768
rect 313332 461728 313338 461740
rect 395522 461728 395528 461740
rect 395580 461728 395586 461780
rect 207198 461660 207204 461712
rect 207256 461700 207262 461712
rect 222838 461700 222844 461712
rect 207256 461672 222844 461700
rect 207256 461660 207262 461672
rect 222838 461660 222844 461672
rect 222896 461660 222902 461712
rect 265066 461660 265072 461712
rect 265124 461700 265130 461712
rect 414658 461700 414664 461712
rect 265124 461672 414664 461700
rect 265124 461660 265130 461672
rect 414658 461660 414664 461672
rect 414716 461660 414722 461712
rect 215478 461592 215484 461644
rect 215536 461632 215542 461644
rect 234614 461632 234620 461644
rect 215536 461604 234620 461632
rect 215536 461592 215542 461604
rect 234614 461592 234620 461604
rect 234672 461592 234678 461644
rect 245654 461592 245660 461644
rect 245712 461632 245718 461644
rect 246390 461632 246396 461644
rect 245712 461604 246396 461632
rect 245712 461592 245718 461604
rect 246390 461592 246396 461604
rect 246448 461592 246454 461644
rect 263778 461592 263784 461644
rect 263836 461632 263842 461644
rect 442994 461632 443000 461644
rect 263836 461604 443000 461632
rect 263836 461592 263842 461604
rect 442994 461592 443000 461604
rect 443052 461592 443058 461644
rect 334066 461524 334072 461576
rect 334124 461564 334130 461576
rect 400766 461564 400772 461576
rect 334124 461536 400772 461564
rect 334124 461524 334130 461536
rect 400766 461524 400772 461536
rect 400824 461524 400830 461576
rect 177482 461456 177488 461508
rect 177540 461496 177546 461508
rect 347774 461496 347780 461508
rect 177540 461468 347780 461496
rect 177540 461456 177546 461468
rect 347774 461456 347780 461468
rect 347832 461456 347838 461508
rect 174814 461388 174820 461440
rect 174872 461428 174878 461440
rect 357434 461428 357440 461440
rect 174872 461400 357440 461428
rect 174872 461388 174878 461400
rect 357434 461388 357440 461400
rect 357492 461388 357498 461440
rect 174906 461320 174912 461372
rect 174964 461360 174970 461372
rect 362954 461360 362960 461372
rect 174964 461332 362960 461360
rect 174964 461320 174970 461332
rect 362954 461320 362960 461332
rect 363012 461320 363018 461372
rect 174722 461252 174728 461304
rect 174780 461292 174786 461304
rect 368474 461292 368480 461304
rect 174780 461264 368480 461292
rect 174780 461252 174786 461264
rect 368474 461252 368480 461264
rect 368532 461252 368538 461304
rect 204438 461184 204444 461236
rect 204496 461224 204502 461236
rect 559558 461224 559564 461236
rect 204496 461196 559564 461224
rect 204496 461184 204502 461196
rect 559558 461184 559564 461196
rect 559616 461184 559622 461236
rect 202874 461116 202880 461168
rect 202932 461156 202938 461168
rect 558270 461156 558276 461168
rect 202932 461128 558276 461156
rect 202932 461116 202938 461128
rect 558270 461116 558276 461128
rect 558328 461116 558334 461168
rect 201494 461048 201500 461100
rect 201552 461088 201558 461100
rect 563698 461088 563704 461100
rect 201552 461060 563704 461088
rect 201552 461048 201558 461060
rect 563698 461048 563704 461060
rect 563756 461048 563762 461100
rect 202966 460980 202972 461032
rect 203024 461020 203030 461032
rect 576118 461020 576124 461032
rect 203024 460992 576124 461020
rect 203024 460980 203030 460992
rect 576118 460980 576124 460992
rect 576176 460980 576182 461032
rect 203058 460912 203064 460964
rect 203116 460952 203122 460964
rect 580718 460952 580724 460964
rect 203116 460924 580724 460952
rect 203116 460912 203122 460924
rect 580718 460912 580724 460924
rect 580776 460912 580782 460964
rect 237558 460776 237564 460828
rect 237616 460816 237622 460828
rect 237926 460816 237932 460828
rect 237616 460788 237932 460816
rect 237616 460776 237622 460788
rect 237926 460776 237932 460788
rect 237984 460776 237990 460828
rect 177390 460572 177396 460624
rect 177448 460612 177454 460624
rect 354858 460612 354864 460624
rect 177448 460584 354864 460612
rect 177448 460572 177454 460584
rect 354858 460572 354864 460584
rect 354916 460572 354922 460624
rect 169294 460504 169300 460556
rect 169352 460544 169358 460556
rect 280982 460544 280988 460556
rect 169352 460516 280988 460544
rect 169352 460504 169358 460516
rect 280982 460504 280988 460516
rect 281040 460504 281046 460556
rect 167822 460436 167828 460488
rect 167880 460476 167886 460488
rect 231302 460476 231308 460488
rect 167880 460448 231308 460476
rect 167880 460436 167886 460448
rect 231302 460436 231308 460448
rect 231360 460436 231366 460488
rect 264422 460436 264428 460488
rect 264480 460476 264486 460488
rect 295978 460476 295984 460488
rect 264480 460448 295984 460476
rect 264480 460436 264486 460448
rect 295978 460436 295984 460448
rect 296036 460436 296042 460488
rect 316126 460436 316132 460488
rect 316184 460476 316190 460488
rect 405366 460476 405372 460488
rect 316184 460448 405372 460476
rect 316184 460436 316190 460448
rect 405366 460436 405372 460448
rect 405424 460436 405430 460488
rect 172054 460368 172060 460420
rect 172112 460408 172118 460420
rect 297542 460408 297548 460420
rect 172112 460380 297548 460408
rect 172112 460368 172118 460380
rect 297542 460368 297548 460380
rect 297600 460368 297606 460420
rect 318794 460368 318800 460420
rect 318852 460408 318858 460420
rect 411806 460408 411812 460420
rect 318852 460380 411812 460408
rect 318852 460368 318858 460380
rect 411806 460368 411812 460380
rect 411864 460368 411870 460420
rect 171962 460300 171968 460352
rect 172020 460340 172026 460352
rect 301590 460340 301596 460352
rect 172020 460312 301596 460340
rect 172020 460300 172026 460312
rect 301590 460300 301596 460312
rect 301648 460300 301654 460352
rect 309226 460300 309232 460352
rect 309284 460340 309290 460352
rect 405274 460340 405280 460352
rect 309284 460312 405280 460340
rect 309284 460300 309290 460312
rect 405274 460300 405280 460312
rect 405332 460300 405338 460352
rect 198366 460232 198372 460284
rect 198424 460272 198430 460284
rect 254486 460272 254492 460284
rect 198424 460244 254492 460272
rect 198424 460232 198430 460244
rect 254486 460232 254492 460244
rect 254544 460232 254550 460284
rect 272150 460232 272156 460284
rect 272208 460272 272214 460284
rect 451274 460272 451280 460284
rect 272208 460244 451280 460272
rect 272208 460232 272214 460244
rect 451274 460232 451280 460244
rect 451332 460232 451338 460284
rect 275462 460164 275468 460216
rect 275520 460204 275526 460216
rect 476758 460204 476764 460216
rect 275520 460176 476764 460204
rect 275520 460164 275526 460176
rect 476758 460164 476764 460176
rect 476816 460164 476822 460216
rect 301038 460096 301044 460148
rect 301096 460136 301102 460148
rect 402514 460136 402520 460148
rect 301096 460108 402520 460136
rect 301096 460096 301102 460108
rect 402514 460096 402520 460108
rect 402572 460096 402578 460148
rect 177666 460028 177672 460080
rect 177724 460068 177730 460080
rect 345750 460068 345756 460080
rect 177724 460040 345756 460068
rect 177724 460028 177730 460040
rect 345750 460028 345756 460040
rect 345808 460028 345814 460080
rect 356790 460028 356796 460080
rect 356848 460068 356854 460080
rect 400950 460068 400956 460080
rect 356848 460040 400956 460068
rect 356848 460028 356854 460040
rect 400950 460028 400956 460040
rect 401008 460028 401014 460080
rect 164142 459960 164148 460012
rect 164200 460000 164206 460012
rect 338390 460000 338396 460012
rect 164200 459972 338396 460000
rect 164200 459960 164206 459972
rect 338390 459960 338396 459972
rect 338448 460000 338454 460012
rect 396718 460000 396724 460012
rect 338448 459972 396724 460000
rect 338448 459960 338454 459972
rect 396718 459960 396724 459972
rect 396776 459960 396782 460012
rect 171870 459892 171876 459944
rect 171928 459932 171934 459944
rect 305638 459932 305644 459944
rect 171928 459904 305644 459932
rect 171928 459892 171934 459904
rect 305638 459892 305644 459904
rect 305696 459892 305702 459944
rect 350902 459892 350908 459944
rect 350960 459932 350966 459944
rect 401042 459932 401048 459944
rect 350960 459904 401048 459932
rect 350960 459892 350966 459904
rect 401042 459892 401048 459904
rect 401100 459892 401106 459944
rect 14918 459824 14924 459876
rect 14976 459864 14982 459876
rect 230566 459864 230572 459876
rect 14976 459836 230572 459864
rect 14976 459824 14982 459836
rect 230566 459824 230572 459836
rect 230624 459824 230630 459876
rect 292758 459824 292764 459876
rect 292816 459864 292822 459876
rect 402238 459864 402244 459876
rect 292816 459836 402244 459864
rect 292816 459824 292822 459836
rect 402238 459824 402244 459836
rect 402296 459824 402302 459876
rect 14458 459756 14464 459808
rect 14516 459796 14522 459808
rect 233326 459796 233332 459808
rect 14516 459768 233332 459796
rect 14516 459756 14522 459768
rect 233326 459756 233332 459768
rect 233384 459756 233390 459808
rect 286502 459756 286508 459808
rect 286560 459796 286566 459808
rect 418890 459796 418896 459808
rect 286560 459768 418896 459796
rect 286560 459756 286566 459768
rect 418890 459756 418896 459768
rect 418948 459756 418954 459808
rect 159818 459688 159824 459740
rect 159876 459728 159882 459740
rect 385494 459728 385500 459740
rect 159876 459700 385500 459728
rect 159876 459688 159882 459700
rect 385494 459688 385500 459700
rect 385552 459688 385558 459740
rect 156690 459620 156696 459672
rect 156748 459660 156754 459672
rect 382550 459660 382556 459672
rect 156748 459632 382556 459660
rect 156748 459620 156754 459632
rect 382550 459620 382556 459632
rect 382608 459620 382614 459672
rect 204530 459552 204536 459604
rect 204588 459592 204594 459604
rect 493410 459592 493416 459604
rect 204588 459564 493416 459592
rect 204588 459552 204594 459564
rect 493410 459552 493416 459564
rect 493468 459552 493474 459604
rect 240134 459484 240140 459536
rect 240192 459524 240198 459536
rect 240870 459524 240876 459536
rect 240192 459496 240876 459524
rect 240192 459484 240198 459496
rect 240870 459484 240876 459496
rect 240928 459484 240934 459536
rect 185670 459280 185676 459332
rect 185728 459320 185734 459332
rect 336182 459320 336188 459332
rect 185728 459292 336188 459320
rect 185728 459280 185734 459292
rect 336182 459280 336188 459292
rect 336240 459280 336246 459332
rect 188522 459212 188528 459264
rect 188580 459252 188586 459264
rect 319622 459252 319628 459264
rect 188580 459224 319628 459252
rect 188580 459212 188586 459224
rect 319622 459212 319628 459224
rect 319680 459212 319686 459264
rect 162486 459144 162492 459196
rect 162544 459184 162550 459196
rect 328546 459184 328552 459196
rect 162544 459156 328552 459184
rect 162544 459144 162550 459156
rect 328546 459144 328552 459156
rect 328604 459144 328610 459196
rect 198182 459076 198188 459128
rect 198240 459116 198246 459128
rect 237374 459116 237380 459128
rect 198240 459088 237380 459116
rect 198240 459076 198246 459088
rect 237374 459076 237380 459088
rect 237432 459076 237438 459128
rect 283650 459076 283656 459128
rect 283708 459116 283714 459128
rect 400858 459116 400864 459128
rect 283708 459088 400864 459116
rect 283708 459076 283714 459088
rect 400858 459076 400864 459088
rect 400916 459076 400922 459128
rect 198090 459008 198096 459060
rect 198148 459048 198154 459060
rect 251358 459048 251364 459060
rect 198148 459020 251364 459048
rect 198148 459008 198154 459020
rect 251358 459008 251364 459020
rect 251416 459008 251422 459060
rect 353846 459008 353852 459060
rect 353904 459048 353910 459060
rect 401134 459048 401140 459060
rect 353904 459020 401140 459048
rect 353904 459008 353910 459020
rect 401134 459008 401140 459020
rect 401192 459008 401198 459060
rect 197998 458940 198004 458992
rect 198056 458980 198062 458992
rect 258074 458980 258080 458992
rect 198056 458952 258080 458980
rect 198056 458940 198062 458952
rect 258074 458940 258080 458952
rect 258132 458940 258138 458992
rect 347958 458940 347964 458992
rect 348016 458980 348022 458992
rect 401226 458980 401232 458992
rect 348016 458952 401232 458980
rect 348016 458940 348022 458952
rect 401226 458940 401232 458952
rect 401284 458940 401290 458992
rect 188890 458872 188896 458924
rect 188948 458912 188954 458924
rect 299658 458912 299664 458924
rect 188948 458884 299664 458912
rect 188948 458872 188954 458884
rect 299658 458872 299664 458884
rect 299716 458872 299722 458924
rect 305178 458872 305184 458924
rect 305236 458912 305242 458924
rect 402422 458912 402428 458924
rect 305236 458884 402428 458912
rect 305236 458872 305242 458884
rect 402422 458872 402428 458884
rect 402480 458872 402486 458924
rect 197354 458804 197360 458856
rect 197412 458844 197418 458856
rect 197538 458844 197544 458856
rect 197412 458816 197544 458844
rect 197412 458804 197418 458816
rect 197538 458804 197544 458816
rect 197596 458804 197602 458856
rect 198274 458804 198280 458856
rect 198332 458844 198338 458856
rect 259454 458844 259460 458856
rect 198332 458816 259460 458844
rect 198332 458804 198338 458816
rect 259454 458804 259460 458816
rect 259512 458804 259518 458856
rect 265526 458804 265532 458856
rect 265584 458844 265590 458856
rect 444374 458844 444380 458856
rect 265584 458816 444380 458844
rect 265584 458804 265590 458816
rect 444374 458804 444380 458816
rect 444432 458804 444438 458856
rect 252830 458736 252836 458788
rect 252888 458776 252894 458788
rect 253014 458776 253020 458788
rect 252888 458748 253020 458776
rect 252888 458736 252894 458748
rect 253014 458736 253020 458748
rect 253072 458736 253078 458788
rect 287974 458736 287980 458788
rect 288032 458776 288038 458788
rect 402330 458776 402336 458788
rect 288032 458748 402336 458776
rect 288032 458736 288038 458748
rect 402330 458736 402336 458748
rect 402388 458736 402394 458788
rect 220998 458668 221004 458720
rect 221056 458708 221062 458720
rect 221366 458708 221372 458720
rect 221056 458680 221372 458708
rect 221056 458668 221062 458680
rect 221366 458668 221372 458680
rect 221424 458668 221430 458720
rect 296806 458668 296812 458720
rect 296864 458708 296870 458720
rect 402606 458708 402612 458720
rect 296864 458680 402612 458708
rect 296864 458668 296870 458680
rect 402606 458668 402612 458680
rect 402664 458668 402670 458720
rect 216766 458600 216772 458652
rect 216824 458640 216830 458652
rect 217686 458640 217692 458652
rect 216824 458612 217692 458640
rect 216824 458600 216830 458612
rect 217686 458600 217692 458612
rect 217744 458600 217750 458652
rect 219526 458600 219532 458652
rect 219584 458640 219590 458652
rect 220262 458640 220268 458652
rect 219584 458612 220268 458640
rect 219584 458600 219590 458612
rect 220262 458600 220268 458612
rect 220320 458600 220326 458652
rect 312630 458600 312636 458652
rect 312688 458640 312694 458652
rect 405458 458640 405464 458652
rect 312688 458612 405464 458640
rect 312688 458600 312694 458612
rect 405458 458600 405464 458612
rect 405516 458600 405522 458652
rect 188614 458532 188620 458584
rect 188672 458572 188678 458584
rect 323118 458572 323124 458584
rect 188672 458544 323124 458572
rect 188672 458532 188678 458544
rect 323118 458532 323124 458544
rect 323176 458532 323182 458584
rect 325694 458532 325700 458584
rect 325752 458572 325758 458584
rect 403986 458572 403992 458584
rect 325752 458544 403992 458572
rect 325752 458532 325758 458544
rect 403986 458532 403992 458544
rect 404044 458532 404050 458584
rect 188338 458464 188344 458516
rect 188396 458504 188402 458516
rect 329926 458504 329932 458516
rect 188396 458476 329932 458504
rect 188396 458464 188402 458476
rect 329926 458464 329932 458476
rect 329984 458464 329990 458516
rect 332686 458464 332692 458516
rect 332744 458504 332750 458516
rect 415302 458504 415308 458516
rect 332744 458476 415308 458504
rect 332744 458464 332750 458476
rect 415302 458464 415308 458476
rect 415360 458464 415366 458516
rect 186958 458396 186964 458448
rect 187016 458436 187022 458448
rect 291194 458436 291200 458448
rect 187016 458408 291200 458436
rect 187016 458396 187022 458408
rect 291194 458396 291200 458408
rect 291252 458396 291258 458448
rect 329190 458396 329196 458448
rect 329248 458436 329254 458448
rect 403894 458436 403900 458448
rect 329248 458408 403900 458436
rect 329248 458396 329254 458408
rect 403894 458396 403900 458408
rect 403952 458396 403958 458448
rect 177574 458328 177580 458380
rect 177632 458368 177638 458380
rect 339862 458368 339868 458380
rect 177632 458340 339868 458368
rect 177632 458328 177638 458340
rect 339862 458328 339868 458340
rect 339920 458328 339926 458380
rect 342438 458328 342444 458380
rect 342496 458368 342502 458380
rect 404078 458368 404084 458380
rect 342496 458340 404084 458368
rect 342496 458328 342502 458340
rect 404078 458328 404084 458340
rect 404136 458328 404142 458380
rect 187050 458260 187056 458312
rect 187108 458300 187114 458312
rect 303982 458300 303988 458312
rect 187108 458272 303988 458300
rect 187108 458260 187114 458272
rect 303982 458260 303988 458272
rect 304040 458260 304046 458312
rect 319254 458260 319260 458312
rect 319312 458300 319318 458312
rect 418798 458300 418804 458312
rect 319312 458272 418804 458300
rect 319312 458260 319318 458272
rect 418798 458260 418804 458272
rect 418856 458260 418862 458312
rect 15010 458192 15016 458244
rect 15068 458232 15074 458244
rect 230658 458232 230664 458244
rect 15068 458204 230664 458232
rect 15068 458192 15074 458204
rect 230658 458192 230664 458204
rect 230716 458192 230722 458244
rect 369946 458192 369952 458244
rect 370004 458232 370010 458244
rect 413370 458232 413376 458244
rect 370004 458204 413376 458232
rect 370004 458192 370010 458204
rect 413370 458192 413376 458204
rect 413428 458192 413434 458244
rect 493410 458124 493416 458176
rect 493468 458164 493474 458176
rect 580166 458164 580172 458176
rect 493468 458136 580172 458164
rect 493468 458124 493474 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 180610 457852 180616 457904
rect 180668 457892 180674 457904
rect 326614 457892 326620 457904
rect 180668 457864 326620 457892
rect 180668 457852 180674 457864
rect 326614 457852 326620 457864
rect 326672 457852 326678 457904
rect 162394 457784 162400 457836
rect 162452 457824 162458 457836
rect 361942 457824 361948 457836
rect 162452 457796 361948 457824
rect 162452 457784 162458 457796
rect 361942 457784 361948 457796
rect 362000 457784 362006 457836
rect 162762 457716 162768 457768
rect 162820 457756 162826 457768
rect 358998 457756 359004 457768
rect 162820 457728 359004 457756
rect 162820 457716 162826 457728
rect 358998 457716 359004 457728
rect 359056 457716 359062 457768
rect 180426 457648 180432 457700
rect 180484 457688 180490 457700
rect 333238 457688 333244 457700
rect 180484 457660 333244 457688
rect 180484 457648 180490 457660
rect 333238 457648 333244 457660
rect 333296 457648 333302 457700
rect 356422 457648 356428 457700
rect 356480 457688 356486 457700
rect 412358 457688 412364 457700
rect 356480 457660 412364 457688
rect 356480 457648 356486 457660
rect 412358 457648 412364 457660
rect 412416 457648 412422 457700
rect 183278 457580 183284 457632
rect 183336 457620 183342 457632
rect 288434 457620 288440 457632
rect 183336 457592 288440 457620
rect 183336 457580 183342 457592
rect 288434 457580 288440 457592
rect 288492 457580 288498 457632
rect 289262 457580 289268 457632
rect 289320 457620 289326 457632
rect 354214 457620 354220 457632
rect 289320 457592 354220 457620
rect 289320 457580 289326 457592
rect 354214 457580 354220 457592
rect 354272 457580 354278 457632
rect 372706 457580 372712 457632
rect 372764 457620 372770 457632
rect 416130 457620 416136 457632
rect 372764 457592 416136 457620
rect 372764 457580 372770 457592
rect 416130 457580 416136 457592
rect 416188 457580 416194 457632
rect 180334 457512 180340 457564
rect 180392 457552 180398 457564
rect 292850 457552 292856 457564
rect 180392 457524 292856 457552
rect 180392 457512 180398 457524
rect 292850 457512 292856 457524
rect 292908 457512 292914 457564
rect 359366 457512 359372 457564
rect 359424 457552 359430 457564
rect 411990 457552 411996 457564
rect 359424 457524 411996 457552
rect 359424 457512 359430 457524
rect 411990 457512 411996 457524
rect 412048 457512 412054 457564
rect 170490 457444 170496 457496
rect 170548 457484 170554 457496
rect 234982 457484 234988 457496
rect 170548 457456 234988 457484
rect 170548 457444 170554 457456
rect 234982 457444 234988 457456
rect 235040 457444 235046 457496
rect 265250 457444 265256 457496
rect 265308 457484 265314 457496
rect 440234 457484 440240 457496
rect 265308 457456 440240 457484
rect 265308 457444 265314 457456
rect 440234 457444 440240 457456
rect 440292 457444 440298 457496
rect 180242 457376 180248 457428
rect 180300 457416 180306 457428
rect 297174 457416 297180 457428
rect 180300 457388 297180 457416
rect 180300 457376 180306 457388
rect 297174 457376 297180 457388
rect 297232 457376 297238 457428
rect 338758 457376 338764 457428
rect 338816 457416 338822 457428
rect 412450 457416 412456 457428
rect 338816 457388 412456 457416
rect 338816 457376 338822 457388
rect 412450 457376 412456 457388
rect 412508 457376 412514 457428
rect 180150 457308 180156 457360
rect 180208 457348 180214 457360
rect 301222 457348 301228 457360
rect 180208 457320 301228 457348
rect 180208 457308 180214 457320
rect 301222 457308 301228 457320
rect 301280 457308 301286 457360
rect 335446 457308 335452 457360
rect 335504 457348 335510 457360
rect 412266 457348 412272 457360
rect 335504 457320 412272 457348
rect 335504 457308 335510 457320
rect 412266 457308 412272 457320
rect 412324 457308 412330 457360
rect 318978 457240 318984 457292
rect 319036 457280 319042 457292
rect 414658 457280 414664 457292
rect 319036 457252 414664 457280
rect 319036 457240 319042 457252
rect 414658 457240 414664 457252
rect 414716 457240 414722 457292
rect 278682 457172 278688 457224
rect 278740 457212 278746 457224
rect 419258 457212 419264 457224
rect 278740 457184 419264 457212
rect 278740 457172 278746 457184
rect 419258 457172 419264 457184
rect 419316 457172 419322 457224
rect 325970 457104 325976 457156
rect 326028 457144 326034 457156
rect 414750 457144 414756 457156
rect 326028 457116 414756 457144
rect 326028 457104 326034 457116
rect 414750 457104 414756 457116
rect 414808 457104 414814 457156
rect 308582 457036 308588 457088
rect 308640 457076 308646 457088
rect 406562 457076 406568 457088
rect 308640 457048 406568 457076
rect 308640 457036 308646 457048
rect 406562 457036 406568 457048
rect 406620 457036 406626 457088
rect 180518 456968 180524 457020
rect 180576 457008 180582 457020
rect 320174 457008 320180 457020
rect 180576 456980 320180 457008
rect 180576 456968 180582 456980
rect 320174 456968 320180 456980
rect 320232 456968 320238 457020
rect 332134 456968 332140 457020
rect 332192 457008 332198 457020
rect 414842 457008 414848 457020
rect 332192 456980 414848 457008
rect 332192 456968 332198 456980
rect 414842 456968 414848 456980
rect 414900 456968 414906 457020
rect 169386 456900 169392 456952
rect 169444 456940 169450 456952
rect 316678 456940 316684 456952
rect 169444 456912 316684 456940
rect 169444 456900 169450 456912
rect 316678 456900 316684 456912
rect 316736 456900 316742 456952
rect 341702 456900 341708 456952
rect 341760 456940 341766 456952
rect 412082 456940 412088 456952
rect 341760 456912 412088 456940
rect 341760 456900 341766 456912
rect 412082 456900 412088 456912
rect 412140 456900 412146 456952
rect 172146 456832 172152 456884
rect 172204 456872 172210 456884
rect 288710 456872 288716 456884
rect 172204 456844 288716 456872
rect 172204 456832 172210 456844
rect 288710 456832 288716 456844
rect 288768 456832 288774 456884
rect 348050 456832 348056 456884
rect 348108 456872 348114 456884
rect 412174 456872 412180 456884
rect 348108 456844 412180 456872
rect 348108 456832 348114 456844
rect 412174 456832 412180 456844
rect 412232 456832 412238 456884
rect 162302 456764 162308 456816
rect 162360 456804 162366 456816
rect 364886 456804 364892 456816
rect 162360 456776 364892 456804
rect 162360 456764 162366 456776
rect 364886 456764 364892 456776
rect 364944 456764 364950 456816
rect 375282 456764 375288 456816
rect 375340 456804 375346 456816
rect 388898 456804 388904 456816
rect 375340 456776 388904 456804
rect 375340 456764 375346 456776
rect 388898 456764 388904 456776
rect 388956 456764 388962 456816
rect 162670 456560 162676 456612
rect 162728 456600 162734 456612
rect 370774 456600 370780 456612
rect 162728 456572 370780 456600
rect 162728 456560 162734 456572
rect 370774 456560 370780 456572
rect 370832 456560 370838 456612
rect 216674 456492 216680 456544
rect 216732 456532 216738 456544
rect 216950 456532 216956 456544
rect 216732 456504 216956 456532
rect 216732 456492 216738 456504
rect 216950 456492 216956 456504
rect 217008 456492 217014 456544
rect 219434 456492 219440 456544
rect 219492 456532 219498 456544
rect 219710 456532 219716 456544
rect 219492 456504 219716 456532
rect 219492 456492 219498 456504
rect 219710 456492 219716 456504
rect 219768 456492 219774 456544
rect 244274 456492 244280 456544
rect 244332 456532 244338 456544
rect 244642 456532 244648 456544
rect 244332 456504 244648 456532
rect 244332 456492 244338 456504
rect 244642 456492 244648 456504
rect 244700 456492 244706 456544
rect 328546 456492 328552 456544
rect 328604 456532 328610 456544
rect 414566 456532 414572 456544
rect 328604 456504 414572 456532
rect 328604 456492 328610 456504
rect 414566 456492 414572 456504
rect 414624 456492 414630 456544
rect 165154 456424 165160 456476
rect 165212 456464 165218 456476
rect 374086 456464 374092 456476
rect 165212 456436 374092 456464
rect 165212 456424 165218 456436
rect 374086 456424 374092 456436
rect 374144 456424 374150 456476
rect 162578 456356 162584 456408
rect 162636 456396 162642 456408
rect 367830 456396 367836 456408
rect 162636 456368 367836 456396
rect 162636 456356 162642 456368
rect 367830 456356 367836 456368
rect 367888 456356 367894 456408
rect 172238 456288 172244 456340
rect 172296 456328 172302 456340
rect 293402 456328 293408 456340
rect 172296 456300 293408 456328
rect 172296 456288 172302 456300
rect 293402 456288 293408 456300
rect 293460 456288 293466 456340
rect 333974 456288 333980 456340
rect 334032 456328 334038 456340
rect 334342 456328 334348 456340
rect 334032 456300 334348 456328
rect 334032 456288 334038 456300
rect 334342 456288 334348 456300
rect 334400 456288 334406 456340
rect 377030 456288 377036 456340
rect 377088 456328 377094 456340
rect 409322 456328 409328 456340
rect 377088 456300 409328 456328
rect 377088 456288 377094 456300
rect 409322 456288 409328 456300
rect 409380 456288 409386 456340
rect 167638 456220 167644 456272
rect 167696 456260 167702 456272
rect 234246 456260 234252 456272
rect 167696 456232 234252 456260
rect 167696 456220 167702 456232
rect 234246 456220 234252 456232
rect 234304 456220 234310 456272
rect 276014 456220 276020 456272
rect 276072 456260 276078 456272
rect 276934 456260 276940 456272
rect 276072 456232 276940 456260
rect 276072 456220 276078 456232
rect 276934 456220 276940 456232
rect 276992 456220 276998 456272
rect 282178 456220 282184 456272
rect 282236 456260 282242 456272
rect 416314 456260 416320 456272
rect 282236 456232 416320 456260
rect 282236 456220 282242 456232
rect 416314 456220 416320 456232
rect 416372 456220 416378 456272
rect 188798 456152 188804 456204
rect 188856 456192 188862 456204
rect 279510 456192 279516 456204
rect 188856 456164 279516 456192
rect 188856 456152 188862 456164
rect 279510 456152 279516 456164
rect 279568 456152 279574 456204
rect 282454 456152 282460 456204
rect 282512 456192 282518 456204
rect 419350 456192 419356 456204
rect 282512 456164 419356 456192
rect 282512 456152 282518 456164
rect 419350 456152 419356 456164
rect 419408 456152 419414 456204
rect 200758 456084 200764 456136
rect 200816 456124 200822 456136
rect 331214 456124 331220 456136
rect 200816 456096 331220 456124
rect 200816 456084 200822 456096
rect 331214 456084 331220 456096
rect 331272 456084 331278 456136
rect 336734 456084 336740 456136
rect 336792 456124 336798 456136
rect 337654 456124 337660 456136
rect 336792 456096 337660 456124
rect 336792 456084 336798 456096
rect 337654 456084 337660 456096
rect 337712 456084 337718 456136
rect 354674 456084 354680 456136
rect 354732 456124 354738 456136
rect 355686 456124 355692 456136
rect 354732 456096 355692 456124
rect 354732 456084 354738 456096
rect 355686 456084 355692 456096
rect 355744 456084 355750 456136
rect 375374 456084 375380 456136
rect 375432 456124 375438 456136
rect 376294 456124 376300 456136
rect 375432 456096 376300 456124
rect 375432 456084 375438 456096
rect 376294 456084 376300 456096
rect 376352 456084 376358 456136
rect 376386 456084 376392 456136
rect 376444 456124 376450 456136
rect 398098 456124 398104 456136
rect 376444 456096 398104 456124
rect 376444 456084 376450 456096
rect 398098 456084 398104 456096
rect 398156 456084 398162 456136
rect 165062 456016 165068 456068
rect 165120 456056 165126 456068
rect 311434 456056 311440 456068
rect 165120 456028 311440 456056
rect 165120 456016 165126 456028
rect 311434 456016 311440 456028
rect 311492 456016 311498 456068
rect 352374 456016 352380 456068
rect 352432 456056 352438 456068
rect 395614 456056 395620 456068
rect 352432 456028 395620 456056
rect 352432 456016 352438 456028
rect 395614 456016 395620 456028
rect 395672 456016 395678 456068
rect 215294 455948 215300 456000
rect 215352 455988 215358 456000
rect 216214 455988 216220 456000
rect 215352 455960 216220 455988
rect 215352 455948 215358 455960
rect 216214 455948 216220 455960
rect 216272 455948 216278 456000
rect 218146 455948 218152 456000
rect 218204 455988 218210 456000
rect 218790 455988 218796 456000
rect 218204 455960 218796 455988
rect 218204 455948 218210 455960
rect 218790 455948 218796 455960
rect 218848 455948 218854 456000
rect 220814 455948 220820 456000
rect 220872 455988 220878 456000
rect 221734 455988 221740 456000
rect 220872 455960 221740 455988
rect 220872 455948 220878 455960
rect 221734 455948 221740 455960
rect 221792 455948 221798 456000
rect 222378 455948 222384 456000
rect 222436 455988 222442 456000
rect 223206 455988 223212 456000
rect 222436 455960 223212 455988
rect 222436 455948 222442 455960
rect 223206 455948 223212 455960
rect 223264 455948 223270 456000
rect 223666 455948 223672 456000
rect 223724 455988 223730 456000
rect 224310 455988 224316 456000
rect 223724 455960 224316 455988
rect 223724 455948 223730 455960
rect 224310 455948 224316 455960
rect 224368 455948 224374 456000
rect 231946 455948 231952 456000
rect 232004 455988 232010 456000
rect 232774 455988 232780 456000
rect 232004 455960 232780 455988
rect 232004 455948 232010 455960
rect 232774 455948 232780 455960
rect 232832 455948 232838 456000
rect 244366 455948 244372 456000
rect 244424 455988 244430 456000
rect 244918 455988 244924 456000
rect 244424 455960 244924 455988
rect 244424 455948 244430 455960
rect 244918 455948 244924 455960
rect 244976 455948 244982 456000
rect 247218 455948 247224 456000
rect 247276 455988 247282 456000
rect 247862 455988 247868 456000
rect 247276 455960 247868 455988
rect 247276 455948 247282 455960
rect 247862 455948 247868 455960
rect 247920 455948 247926 456000
rect 251174 455948 251180 456000
rect 251232 455988 251238 456000
rect 251910 455988 251916 456000
rect 251232 455960 251916 455988
rect 251232 455948 251238 455960
rect 251910 455948 251916 455960
rect 251968 455948 251974 456000
rect 252646 455948 252652 456000
rect 252704 455988 252710 456000
rect 253382 455988 253388 456000
rect 252704 455960 253388 455988
rect 252704 455948 252710 455960
rect 253382 455948 253388 455960
rect 253440 455948 253446 456000
rect 273346 455948 273352 456000
rect 273404 455988 273410 456000
rect 273990 455988 273996 456000
rect 273404 455960 273996 455988
rect 273404 455948 273410 455960
rect 273990 455948 273996 455960
rect 274048 455948 274054 456000
rect 276106 455948 276112 456000
rect 276164 455988 276170 456000
rect 276566 455988 276572 456000
rect 276164 455960 276572 455988
rect 276164 455948 276170 455960
rect 276566 455948 276572 455960
rect 276624 455948 276630 456000
rect 312262 455948 312268 456000
rect 312320 455988 312326 456000
rect 403710 455988 403716 456000
rect 312320 455960 403716 455988
rect 312320 455948 312326 455960
rect 403710 455948 403716 455960
rect 403768 455948 403774 456000
rect 164050 455880 164056 455932
rect 164108 455920 164114 455932
rect 316310 455920 316316 455932
rect 164108 455892 316316 455920
rect 164108 455880 164114 455892
rect 316310 455880 316316 455892
rect 316368 455880 316374 455932
rect 339126 455880 339132 455932
rect 339184 455920 339190 455932
rect 404170 455920 404176 455932
rect 339184 455892 404176 455920
rect 339184 455880 339190 455892
rect 404170 455880 404176 455892
rect 404228 455880 404234 455932
rect 191190 455812 191196 455864
rect 191248 455852 191254 455864
rect 200758 455852 200764 455864
rect 191248 455824 200764 455852
rect 191248 455812 191254 455824
rect 200758 455812 200764 455824
rect 200816 455812 200822 455864
rect 322198 455812 322204 455864
rect 322256 455852 322262 455864
rect 414934 455852 414940 455864
rect 322256 455824 414940 455852
rect 322256 455812 322262 455824
rect 414934 455812 414940 455824
rect 414992 455812 414998 455864
rect 158070 455744 158076 455796
rect 158128 455784 158134 455796
rect 330018 455784 330024 455796
rect 158128 455756 330024 455784
rect 158128 455744 158134 455756
rect 330018 455744 330024 455756
rect 330076 455744 330082 455796
rect 374454 455744 374460 455796
rect 374512 455784 374518 455796
rect 376386 455784 376392 455796
rect 374512 455756 376392 455784
rect 374512 455744 374518 455756
rect 376386 455744 376392 455756
rect 376444 455744 376450 455796
rect 158254 455676 158260 455728
rect 158312 455716 158318 455728
rect 322934 455716 322940 455728
rect 158312 455688 322940 455716
rect 158312 455676 158318 455688
rect 322934 455676 322940 455688
rect 322992 455676 322998 455728
rect 358262 455676 358268 455728
rect 358320 455716 358326 455728
rect 392946 455716 392952 455728
rect 358320 455688 392952 455716
rect 358320 455676 358326 455688
rect 392946 455676 392952 455688
rect 393004 455676 393010 455728
rect 273438 455608 273444 455660
rect 273496 455648 273502 455660
rect 273622 455648 273628 455660
rect 273496 455620 273628 455648
rect 273496 455608 273502 455620
rect 273622 455608 273628 455620
rect 273680 455608 273686 455660
rect 368658 455608 368664 455660
rect 368716 455648 368722 455660
rect 409230 455648 409236 455660
rect 368716 455620 409236 455648
rect 368716 455608 368722 455620
rect 409230 455608 409236 455620
rect 409288 455608 409294 455660
rect 162210 455540 162216 455592
rect 162268 455580 162274 455592
rect 313366 455580 313372 455592
rect 162268 455552 313372 455580
rect 162268 455540 162274 455552
rect 313366 455540 313372 455552
rect 313424 455540 313430 455592
rect 371510 455540 371516 455592
rect 371568 455580 371574 455592
rect 398190 455580 398196 455592
rect 371568 455552 398196 455580
rect 371568 455540 371574 455552
rect 398190 455540 398196 455552
rect 398248 455540 398254 455592
rect 164970 455472 164976 455524
rect 165028 455512 165034 455524
rect 376754 455512 376760 455524
rect 165028 455484 376760 455512
rect 165028 455472 165034 455484
rect 376754 455472 376760 455484
rect 376812 455472 376818 455524
rect 377398 455472 377404 455524
rect 377456 455512 377462 455524
rect 398282 455512 398288 455524
rect 377456 455484 398288 455512
rect 377456 455472 377462 455484
rect 398282 455472 398288 455484
rect 398340 455472 398346 455524
rect 164878 455404 164884 455456
rect 164936 455444 164942 455456
rect 379882 455444 379888 455456
rect 164936 455416 379888 455444
rect 164936 455404 164942 455416
rect 379882 455404 379888 455416
rect 379940 455404 379946 455456
rect 381722 455404 381728 455456
rect 381780 455444 381786 455456
rect 416222 455444 416228 455456
rect 381780 455416 416228 455444
rect 381780 455404 381786 455416
rect 416222 455404 416228 455416
rect 416280 455404 416286 455456
rect 18966 455064 18972 455116
rect 19024 455104 19030 455116
rect 299474 455104 299480 455116
rect 19024 455076 299480 455104
rect 19024 455064 19030 455076
rect 299474 455064 299480 455076
rect 299532 455064 299538 455116
rect 19058 454996 19064 455048
rect 19116 455036 19122 455048
rect 295978 455036 295984 455048
rect 19116 455008 295984 455036
rect 19116 454996 19122 455008
rect 295978 454996 295984 455008
rect 296036 454996 296042 455048
rect 306650 454996 306656 455048
rect 306708 455036 306714 455048
rect 394326 455036 394332 455048
rect 306708 455008 394332 455036
rect 306708 454996 306714 455008
rect 394326 454996 394332 455008
rect 394384 454996 394390 455048
rect 188982 454928 188988 454980
rect 189040 454968 189046 454980
rect 278038 454968 278044 454980
rect 189040 454940 278044 454968
rect 189040 454928 189046 454940
rect 278038 454928 278044 454940
rect 278096 454968 278102 454980
rect 278682 454968 278688 454980
rect 278096 454940 278688 454968
rect 278096 454928 278102 454940
rect 278682 454928 278688 454940
rect 278740 454928 278746 454980
rect 328822 454928 328828 454980
rect 328880 454968 328886 454980
rect 415026 454968 415032 454980
rect 328880 454940 415032 454968
rect 328880 454928 328886 454940
rect 415026 454928 415032 454940
rect 415084 454928 415090 454980
rect 166902 454860 166908 454912
rect 166960 454900 166966 454912
rect 285950 454900 285956 454912
rect 166960 454872 285956 454900
rect 166960 454860 166966 454872
rect 285950 454860 285956 454872
rect 286008 454860 286014 454912
rect 317506 454860 317512 454912
rect 317564 454900 317570 454912
rect 388530 454900 388536 454912
rect 317564 454872 388536 454900
rect 317564 454860 317570 454872
rect 388530 454860 388536 454872
rect 388588 454860 388594 454912
rect 191282 454792 191288 454844
rect 191340 454832 191346 454844
rect 321830 454832 321836 454844
rect 191340 454804 321836 454832
rect 191340 454792 191346 454804
rect 321830 454792 321836 454804
rect 321888 454832 321894 454844
rect 321888 454804 325694 454832
rect 321888 454792 321894 454804
rect 169478 454724 169484 454776
rect 169536 454764 169542 454776
rect 309962 454764 309968 454776
rect 169536 454736 309968 454764
rect 169536 454724 169542 454736
rect 309962 454724 309968 454736
rect 310020 454724 310026 454776
rect 325666 454764 325694 454804
rect 331214 454792 331220 454844
rect 331272 454832 331278 454844
rect 331766 454832 331772 454844
rect 331272 454804 331772 454832
rect 331272 454792 331278 454804
rect 331766 454792 331772 454804
rect 331824 454832 331830 454844
rect 389910 454832 389916 454844
rect 331824 454804 389916 454832
rect 331824 454792 331830 454804
rect 389910 454792 389916 454804
rect 389968 454792 389974 454844
rect 396810 454764 396816 454776
rect 325666 454736 396816 454764
rect 396810 454724 396816 454736
rect 396868 454724 396874 454776
rect 168098 454656 168104 454708
rect 168156 454696 168162 454708
rect 310514 454696 310520 454708
rect 168156 454668 310520 454696
rect 168156 454656 168162 454668
rect 310514 454656 310520 454668
rect 310572 454656 310578 454708
rect 314102 454656 314108 454708
rect 314160 454696 314166 454708
rect 394142 454696 394148 454708
rect 314160 454668 394148 454696
rect 314160 454656 314166 454668
rect 394142 454656 394148 454668
rect 394200 454656 394206 454708
rect 172330 454588 172336 454640
rect 172388 454628 172394 454640
rect 344554 454628 344560 454640
rect 172388 454600 344560 454628
rect 172388 454588 172394 454600
rect 344554 454588 344560 454600
rect 344612 454588 344618 454640
rect 169662 454520 169668 454572
rect 169720 454560 169726 454572
rect 347498 454560 347504 454572
rect 169720 454532 347504 454560
rect 169720 454520 169726 454532
rect 347498 454520 347504 454532
rect 347556 454520 347562 454572
rect 363138 454520 363144 454572
rect 363196 454560 363202 454572
rect 401318 454560 401324 454572
rect 363196 454532 401324 454560
rect 363196 454520 363202 454532
rect 401318 454520 401324 454532
rect 401376 454520 401382 454572
rect 161290 454452 161296 454504
rect 161348 454492 161354 454504
rect 353294 454492 353300 454504
rect 161348 454464 353300 454492
rect 161348 454452 161354 454464
rect 353294 454452 353300 454464
rect 353352 454452 353358 454504
rect 361206 454452 361212 454504
rect 361264 454492 361270 454504
rect 418982 454492 418988 454504
rect 361264 454464 418988 454492
rect 361264 454452 361270 454464
rect 418982 454452 418988 454464
rect 419040 454452 419046 454504
rect 14826 454384 14832 454436
rect 14884 454424 14890 454436
rect 230934 454424 230940 454436
rect 14884 454396 230940 454424
rect 14884 454384 14890 454396
rect 230934 454384 230940 454396
rect 230992 454384 230998 454436
rect 285030 454384 285036 454436
rect 285088 454424 285094 454436
rect 391290 454424 391296 454436
rect 285088 454396 391296 454424
rect 285088 454384 285094 454396
rect 391290 454384 391296 454396
rect 391348 454384 391354 454436
rect 289446 454316 289452 454368
rect 289504 454356 289510 454368
rect 391382 454356 391388 454368
rect 289504 454328 391388 454356
rect 289504 454316 289510 454328
rect 391382 454316 391388 454328
rect 391440 454316 391446 454368
rect 294138 454248 294144 454300
rect 294196 454288 294202 454300
rect 391198 454288 391204 454300
rect 294196 454260 391204 454288
rect 294196 454248 294202 454260
rect 391198 454248 391204 454260
rect 391256 454248 391262 454300
rect 18874 454180 18880 454232
rect 18932 454220 18938 454232
rect 304074 454220 304080 454232
rect 18932 454192 304080 454220
rect 18932 454180 18938 454192
rect 304074 454180 304080 454192
rect 304132 454220 304138 454232
rect 304718 454220 304724 454232
rect 304132 454192 304724 454220
rect 304132 454180 304138 454192
rect 304718 454180 304724 454192
rect 304776 454180 304782 454232
rect 310698 454180 310704 454232
rect 310756 454220 310762 454232
rect 394234 454220 394240 454232
rect 310756 454192 394240 454220
rect 310756 454180 310762 454192
rect 394234 454180 394240 454192
rect 394292 454180 394298 454232
rect 18782 454112 18788 454164
rect 18840 454152 18846 454164
rect 308122 454152 308128 454164
rect 18840 454124 308128 454152
rect 18840 454112 18846 454124
rect 308122 454112 308128 454124
rect 308180 454112 308186 454164
rect 375926 454112 375932 454164
rect 375984 454152 375990 454164
rect 392762 454152 392768 454164
rect 375984 454124 392768 454152
rect 375984 454112 375990 454124
rect 392762 454112 392768 454124
rect 392820 454112 392826 454164
rect 19334 454044 19340 454096
rect 19392 454084 19398 454096
rect 312170 454084 312176 454096
rect 19392 454056 312176 454084
rect 19392 454044 19398 454056
rect 312170 454044 312176 454056
rect 312228 454044 312234 454096
rect 384298 454044 384304 454096
rect 384356 454084 384362 454096
rect 389358 454084 389364 454096
rect 384356 454056 389364 454084
rect 384356 454044 384362 454056
rect 389358 454044 389364 454056
rect 389416 454044 389422 454096
rect 175090 453636 175096 453688
rect 175148 453676 175154 453688
rect 341610 453676 341616 453688
rect 175148 453648 341616 453676
rect 175148 453636 175154 453648
rect 341610 453636 341616 453648
rect 341668 453636 341674 453688
rect 347866 453636 347872 453688
rect 347924 453676 347930 453688
rect 348050 453676 348056 453688
rect 347924 453648 348056 453676
rect 347924 453636 347930 453648
rect 348050 453636 348056 453648
rect 348108 453636 348114 453688
rect 17402 453568 17408 453620
rect 17460 453608 17466 453620
rect 291654 453608 291660 453620
rect 17460 453580 291660 453608
rect 17460 453568 17466 453580
rect 291654 453568 291660 453580
rect 291712 453568 291718 453620
rect 304718 453568 304724 453620
rect 304776 453608 304782 453620
rect 417510 453608 417516 453620
rect 304776 453580 417516 453608
rect 304776 453568 304782 453580
rect 417510 453568 417516 453580
rect 417568 453568 417574 453620
rect 214098 453500 214104 453552
rect 214156 453540 214162 453552
rect 214742 453540 214748 453552
rect 214156 453512 214748 453540
rect 214156 453500 214162 453512
rect 214742 453500 214748 453512
rect 214800 453500 214806 453552
rect 258258 453500 258264 453552
rect 258316 453540 258322 453552
rect 258902 453540 258908 453552
rect 258316 453512 258908 453540
rect 258316 453500 258322 453512
rect 258902 453500 258908 453512
rect 258960 453500 258966 453552
rect 269298 453500 269304 453552
rect 269356 453540 269362 453552
rect 269942 453540 269948 453552
rect 269356 453512 269948 453540
rect 269356 453500 269362 453512
rect 269942 453500 269948 453512
rect 270000 453500 270006 453552
rect 273162 453500 273168 453552
rect 273220 453540 273226 453552
rect 283558 453540 283564 453552
rect 273220 453512 283564 453540
rect 273220 453500 273226 453512
rect 283558 453500 283564 453512
rect 283616 453500 283622 453552
rect 299474 453500 299480 453552
rect 299532 453540 299538 453552
rect 300026 453540 300032 453552
rect 299532 453512 300032 453540
rect 299532 453500 299538 453512
rect 300026 453500 300032 453512
rect 300084 453540 300090 453552
rect 390278 453540 390284 453552
rect 300084 453512 390284 453540
rect 300084 453500 300090 453512
rect 390278 453500 390284 453512
rect 390336 453500 390342 453552
rect 191466 453432 191472 453484
rect 191524 453472 191530 453484
rect 282454 453472 282460 453484
rect 191524 453444 282460 453472
rect 191524 453432 191530 453444
rect 282454 453432 282460 453444
rect 282512 453432 282518 453484
rect 295978 453432 295984 453484
rect 296036 453472 296042 453484
rect 390186 453472 390192 453484
rect 296036 453444 390192 453472
rect 296036 453432 296042 453444
rect 390186 453432 390192 453444
rect 390244 453432 390250 453484
rect 189810 453364 189816 453416
rect 189868 453404 189874 453416
rect 325050 453404 325056 453416
rect 189868 453376 325056 453404
rect 189868 453364 189874 453376
rect 325050 453364 325056 453376
rect 325108 453364 325114 453416
rect 343818 453364 343824 453416
rect 343876 453404 343882 453416
rect 343876 453376 350534 453404
rect 343876 453364 343882 453376
rect 182726 453296 182732 453348
rect 182784 453336 182790 453348
rect 328362 453336 328368 453348
rect 182784 453308 328368 453336
rect 182784 453296 182790 453308
rect 328362 453296 328368 453308
rect 328420 453296 328426 453348
rect 340874 453296 340880 453348
rect 340932 453336 340938 453348
rect 340932 453308 350028 453336
rect 340932 453296 340938 453308
rect 179966 453228 179972 453280
rect 180024 453268 180030 453280
rect 331674 453268 331680 453280
rect 180024 453240 331680 453268
rect 180024 453228 180030 453240
rect 331674 453228 331680 453240
rect 331732 453228 331738 453280
rect 177206 453160 177212 453212
rect 177264 453200 177270 453212
rect 338114 453200 338120 453212
rect 177264 453172 338120 453200
rect 177264 453160 177270 453172
rect 338114 453160 338120 453172
rect 338172 453160 338178 453212
rect 342254 453160 342260 453212
rect 342312 453200 342318 453212
rect 343174 453200 343180 453212
rect 342312 453172 343180 453200
rect 342312 453160 342318 453172
rect 343174 453160 343180 453172
rect 343232 453160 343238 453212
rect 349154 453160 349160 453212
rect 349212 453200 349218 453212
rect 349798 453200 349804 453212
rect 349212 453172 349804 453200
rect 349212 453160 349218 453172
rect 349798 453160 349804 453172
rect 349856 453160 349862 453212
rect 350000 453200 350028 453308
rect 350506 453268 350534 453376
rect 371234 453296 371240 453348
rect 371292 453336 371298 453348
rect 375282 453336 375288 453348
rect 371292 453308 375288 453336
rect 371292 453296 371298 453308
rect 375282 453296 375288 453308
rect 375340 453296 375346 453348
rect 395798 453268 395804 453280
rect 350506 453240 395804 453268
rect 395798 453228 395804 453240
rect 395856 453228 395862 453280
rect 395890 453200 395896 453212
rect 350000 453172 395896 453200
rect 395890 453160 395896 453172
rect 395948 453160 395954 453212
rect 191374 453092 191380 453144
rect 191432 453132 191438 453144
rect 356054 453132 356060 453144
rect 191432 453104 356060 453132
rect 191432 453092 191438 453104
rect 356054 453092 356060 453104
rect 356112 453092 356118 453144
rect 364334 453092 364340 453144
rect 364392 453132 364398 453144
rect 393130 453132 393136 453144
rect 364392 453104 393136 453132
rect 364392 453092 364398 453104
rect 393130 453092 393136 453104
rect 393188 453092 393194 453144
rect 17770 453024 17776 453076
rect 17828 453064 17834 453076
rect 17828 453036 277394 453064
rect 17828 453024 17834 453036
rect 4062 452956 4068 453008
rect 4120 452996 4126 453008
rect 226058 452996 226064 453008
rect 4120 452968 226064 452996
rect 4120 452956 4126 452968
rect 226058 452956 226064 452968
rect 226116 452956 226122 453008
rect 234706 452956 234712 453008
rect 234764 452996 234770 453008
rect 235350 452996 235356 453008
rect 234764 452968 235356 452996
rect 234764 452956 234770 452968
rect 235350 452956 235356 452968
rect 235408 452956 235414 453008
rect 236086 452956 236092 453008
rect 236144 452996 236150 453008
rect 236546 452996 236552 453008
rect 236144 452968 236552 452996
rect 236144 452956 236150 452968
rect 236546 452956 236552 452968
rect 236604 452956 236610 453008
rect 237466 452956 237472 453008
rect 237524 452996 237530 453008
rect 238294 452996 238300 453008
rect 237524 452968 238300 452996
rect 237524 452956 237530 452968
rect 238294 452956 238300 452968
rect 238352 452956 238358 453008
rect 238938 452956 238944 453008
rect 238996 452996 239002 453008
rect 239122 452996 239128 453008
rect 238996 452968 239128 452996
rect 238996 452956 239002 452968
rect 239122 452956 239128 452968
rect 239180 452956 239186 453008
rect 241514 452956 241520 453008
rect 241572 452996 241578 453008
rect 242342 452996 242348 453008
rect 241572 452968 242348 452996
rect 241572 452956 241578 452968
rect 242342 452956 242348 452968
rect 242400 452956 242406 453008
rect 242986 452956 242992 453008
rect 243044 452996 243050 453008
rect 243446 452996 243452 453008
rect 243044 452968 243452 452996
rect 243044 452956 243050 452968
rect 243446 452956 243452 452968
rect 243504 452956 243510 453008
rect 254118 452956 254124 453008
rect 254176 452996 254182 453008
rect 254854 452996 254860 453008
rect 254176 452968 254860 452996
rect 254176 452956 254182 452968
rect 254854 452956 254860 452968
rect 254912 452956 254918 453008
rect 255314 452956 255320 453008
rect 255372 452996 255378 453008
rect 255958 452996 255964 453008
rect 255372 452968 255964 452996
rect 255372 452956 255378 452968
rect 255958 452956 255964 452968
rect 256016 452956 256022 453008
rect 256786 452956 256792 453008
rect 256844 452996 256850 453008
rect 257062 452996 257068 453008
rect 256844 452968 257068 452996
rect 256844 452956 256850 452968
rect 257062 452956 257068 452968
rect 257120 452956 257126 453008
rect 258074 452956 258080 453008
rect 258132 452996 258138 453008
rect 258258 452996 258264 453008
rect 258132 452968 258264 452996
rect 258132 452956 258138 452968
rect 258258 452956 258264 452968
rect 258316 452956 258322 453008
rect 259546 452956 259552 453008
rect 259604 452996 259610 453008
rect 260374 452996 260380 453008
rect 259604 452968 260380 452996
rect 259604 452956 259610 452968
rect 260374 452956 260380 452968
rect 260432 452956 260438 453008
rect 260926 452956 260932 453008
rect 260984 452996 260990 453008
rect 261478 452996 261484 453008
rect 260984 452968 261484 452996
rect 260984 452956 260990 452968
rect 261478 452956 261484 452968
rect 261536 452956 261542 453008
rect 262214 452956 262220 453008
rect 262272 452996 262278 453008
rect 262950 452996 262956 453008
rect 262272 452968 262956 452996
rect 262272 452956 262278 452968
rect 262950 452956 262956 452968
rect 263008 452956 263014 453008
rect 263594 452956 263600 453008
rect 263652 452996 263658 453008
rect 263778 452996 263784 453008
rect 263652 452968 263784 452996
rect 263652 452956 263658 452968
rect 263778 452956 263784 452968
rect 263836 452956 263842 453008
rect 269114 452956 269120 453008
rect 269172 452996 269178 453008
rect 269298 452996 269304 453008
rect 269172 452968 269304 452996
rect 269172 452956 269178 452968
rect 269298 452956 269304 452968
rect 269356 452956 269362 453008
rect 270678 452956 270684 453008
rect 270736 452996 270742 453008
rect 271414 452996 271420 453008
rect 270736 452968 271420 452996
rect 270736 452956 270742 452968
rect 271414 452956 271420 452968
rect 271472 452956 271478 453008
rect 271874 452956 271880 453008
rect 271932 452996 271938 453008
rect 272518 452996 272524 453008
rect 271932 452968 272524 452996
rect 271932 452956 271938 452968
rect 272518 452956 272524 452968
rect 272576 452956 272582 453008
rect 3418 452888 3424 452940
rect 3476 452928 3482 452940
rect 227530 452928 227536 452940
rect 3476 452900 227536 452928
rect 3476 452888 3482 452900
rect 227530 452888 227536 452900
rect 227588 452888 227594 452940
rect 236178 452888 236184 452940
rect 236236 452928 236242 452940
rect 236822 452928 236828 452940
rect 236236 452900 236828 452928
rect 236236 452888 236242 452900
rect 236822 452888 236828 452900
rect 236880 452888 236886 452940
rect 238754 452888 238760 452940
rect 238812 452928 238818 452940
rect 239398 452928 239404 452940
rect 238812 452900 239404 452928
rect 238812 452888 238818 452900
rect 239398 452888 239404 452900
rect 239456 452888 239462 452940
rect 256694 452888 256700 452940
rect 256752 452928 256758 452940
rect 257430 452928 257436 452940
rect 256752 452900 257436 452928
rect 256752 452888 256758 452900
rect 257430 452888 257436 452900
rect 257488 452888 257494 452940
rect 259638 452888 259644 452940
rect 259696 452928 259702 452940
rect 260006 452928 260012 452940
rect 259696 452900 260012 452928
rect 259696 452888 259702 452900
rect 260006 452888 260012 452900
rect 260064 452888 260070 452940
rect 270586 452888 270592 452940
rect 270644 452928 270650 452940
rect 271046 452928 271052 452940
rect 270644 452900 271052 452928
rect 270644 452888 270650 452900
rect 271046 452888 271052 452900
rect 271104 452888 271110 452940
rect 277366 452928 277394 453036
rect 302326 453024 302332 453076
rect 302384 453064 302390 453076
rect 302694 453064 302700 453076
rect 302384 453036 302700 453064
rect 302384 453024 302390 453036
rect 302694 453024 302700 453036
rect 302752 453024 302758 453076
rect 337562 453024 337568 453076
rect 337620 453064 337626 453076
rect 398650 453064 398656 453076
rect 337620 453036 398656 453064
rect 337620 453024 337626 453036
rect 398650 453024 398656 453036
rect 398708 453024 398714 453076
rect 291654 452956 291660 453008
rect 291712 452996 291718 453008
rect 390094 452996 390100 453008
rect 291712 452968 390100 452996
rect 291712 452956 291718 452968
rect 390094 452956 390100 452968
rect 390152 452956 390158 453008
rect 287146 452928 287152 452940
rect 277366 452900 287152 452928
rect 287146 452888 287152 452900
rect 287204 452928 287210 452940
rect 388806 452928 388812 452940
rect 287204 452900 388812 452928
rect 287204 452888 287210 452900
rect 388806 452888 388812 452900
rect 388864 452888 388870 452940
rect 3326 452820 3332 452872
rect 3384 452860 3390 452872
rect 226426 452860 226432 452872
rect 3384 452832 226432 452860
rect 3384 452820 3390 452832
rect 226426 452820 226432 452832
rect 226484 452820 226490 452872
rect 238846 452820 238852 452872
rect 238904 452860 238910 452872
rect 239766 452860 239772 452872
rect 238904 452832 239772 452860
rect 238904 452820 238910 452832
rect 239766 452820 239772 452832
rect 239824 452820 239830 452872
rect 312170 452820 312176 452872
rect 312228 452860 312234 452872
rect 417694 452860 417700 452872
rect 312228 452832 417700 452860
rect 312228 452820 312234 452832
rect 417694 452820 417700 452832
rect 417752 452820 417758 452872
rect 3786 452752 3792 452804
rect 3844 452792 3850 452804
rect 228634 452792 228640 452804
rect 3844 452764 228640 452792
rect 3844 452752 3850 452764
rect 228634 452752 228640 452764
rect 228692 452752 228698 452804
rect 308122 452752 308128 452804
rect 308180 452792 308186 452804
rect 417602 452792 417608 452804
rect 308180 452764 417608 452792
rect 308180 452752 308186 452764
rect 417602 452752 417608 452764
rect 417660 452752 417666 452804
rect 198734 452684 198740 452736
rect 198792 452724 198798 452736
rect 199286 452724 199292 452736
rect 198792 452696 199292 452724
rect 198792 452684 198798 452696
rect 199286 452684 199292 452696
rect 199344 452684 199350 452736
rect 202874 452684 202880 452736
rect 202932 452724 202938 452736
rect 203702 452724 203708 452736
rect 202932 452696 203708 452724
rect 202932 452684 202938 452696
rect 203702 452684 203708 452696
rect 203760 452684 203766 452736
rect 204346 452684 204352 452736
rect 204404 452724 204410 452736
rect 204806 452724 204812 452736
rect 204404 452696 204812 452724
rect 204404 452684 204410 452696
rect 204806 452684 204812 452696
rect 204864 452684 204870 452736
rect 205818 452684 205824 452736
rect 205876 452724 205882 452736
rect 206278 452724 206284 452736
rect 205876 452696 206284 452724
rect 205876 452684 205882 452696
rect 206278 452684 206284 452696
rect 206336 452684 206342 452736
rect 207014 452684 207020 452736
rect 207072 452724 207078 452736
rect 207382 452724 207388 452736
rect 207072 452696 207388 452724
rect 207072 452684 207078 452696
rect 207382 452684 207388 452696
rect 207440 452684 207446 452736
rect 208486 452684 208492 452736
rect 208544 452724 208550 452736
rect 209222 452724 209228 452736
rect 208544 452696 209228 452724
rect 208544 452684 208550 452696
rect 209222 452684 209228 452696
rect 209280 452684 209286 452736
rect 209866 452684 209872 452736
rect 209924 452724 209930 452736
rect 210326 452724 210332 452736
rect 209924 452696 210332 452724
rect 209924 452684 209930 452696
rect 210326 452684 210332 452696
rect 210384 452684 210390 452736
rect 211154 452684 211160 452736
rect 211212 452724 211218 452736
rect 211430 452724 211436 452736
rect 211212 452696 211436 452724
rect 211212 452684 211218 452696
rect 211430 452684 211436 452696
rect 211488 452684 211494 452736
rect 212534 452684 212540 452736
rect 212592 452724 212598 452736
rect 212902 452724 212908 452736
rect 212592 452696 212908 452724
rect 212592 452684 212598 452696
rect 212902 452684 212908 452696
rect 212960 452684 212966 452736
rect 213914 452684 213920 452736
rect 213972 452724 213978 452736
rect 214098 452724 214104 452736
rect 213972 452696 214104 452724
rect 213972 452684 213978 452696
rect 214098 452684 214104 452696
rect 214156 452684 214162 452736
rect 287514 452684 287520 452736
rect 287572 452724 287578 452736
rect 416958 452724 416964 452736
rect 287572 452696 416964 452724
rect 287572 452684 287578 452696
rect 416958 452684 416964 452696
rect 417016 452684 417022 452736
rect 193858 452616 193864 452668
rect 193916 452656 193922 452668
rect 224954 452656 224960 452668
rect 193916 452628 224960 452656
rect 193916 452616 193922 452628
rect 224954 452616 224960 452628
rect 225012 452616 225018 452668
rect 370314 452616 370320 452668
rect 370372 452656 370378 452668
rect 392854 452656 392860 452668
rect 370372 452628 392860 452656
rect 370372 452616 370378 452628
rect 392854 452616 392860 452628
rect 392912 452616 392918 452668
rect 198826 452548 198832 452600
rect 198884 452588 198890 452600
rect 199654 452588 199660 452600
rect 198884 452560 199660 452588
rect 198884 452548 198890 452560
rect 199654 452548 199660 452560
rect 199712 452548 199718 452600
rect 204254 452548 204260 452600
rect 204312 452588 204318 452600
rect 205174 452588 205180 452600
rect 204312 452560 205180 452588
rect 204312 452548 204318 452560
rect 205174 452548 205180 452560
rect 205232 452548 205238 452600
rect 205726 452548 205732 452600
rect 205784 452588 205790 452600
rect 206646 452588 206652 452600
rect 205784 452560 206652 452588
rect 205784 452548 205790 452560
rect 206646 452548 206652 452560
rect 206704 452548 206710 452600
rect 209774 452548 209780 452600
rect 209832 452588 209838 452600
rect 210694 452588 210700 452600
rect 209832 452560 210700 452588
rect 209832 452548 209838 452560
rect 210694 452548 210700 452560
rect 210752 452548 210758 452600
rect 212626 452548 212632 452600
rect 212684 452588 212690 452600
rect 213270 452588 213276 452600
rect 212684 452560 213276 452588
rect 212684 452548 212690 452560
rect 213270 452548 213276 452560
rect 213328 452548 213334 452600
rect 299658 452480 299664 452532
rect 299716 452520 299722 452532
rect 303890 452520 303896 452532
rect 299716 452492 303896 452520
rect 299716 452480 299722 452492
rect 303890 452480 303896 452492
rect 303948 452480 303954 452532
rect 302206 452288 311894 452316
rect 156966 452208 156972 452260
rect 157024 452248 157030 452260
rect 294874 452248 294880 452260
rect 157024 452220 294880 452248
rect 157024 452208 157030 452220
rect 294874 452208 294880 452220
rect 294932 452208 294938 452260
rect 163406 452140 163412 452192
rect 163464 452180 163470 452192
rect 302206 452180 302234 452288
rect 163464 452152 302234 452180
rect 163464 452140 163470 452152
rect 303706 452140 303712 452192
rect 303764 452180 303770 452192
rect 304258 452180 304264 452192
rect 303764 452152 304264 452180
rect 303764 452140 303770 452152
rect 304258 452140 304264 452152
rect 304316 452140 304322 452192
rect 311866 452180 311894 452288
rect 367370 452276 367376 452328
rect 367428 452316 367434 452328
rect 375190 452316 375196 452328
rect 367428 452288 375196 452316
rect 367428 452276 367434 452288
rect 375190 452276 375196 452288
rect 375248 452276 375254 452328
rect 385034 452276 385040 452328
rect 385092 452316 385098 452328
rect 394418 452316 394424 452328
rect 385092 452288 394424 452316
rect 385092 452276 385098 452288
rect 394418 452276 394424 452288
rect 394476 452276 394482 452328
rect 325418 452208 325424 452260
rect 325476 452248 325482 452260
rect 387702 452248 387708 452260
rect 325476 452220 387708 452248
rect 325476 452208 325482 452220
rect 387702 452208 387708 452220
rect 387760 452208 387766 452260
rect 335354 452180 335360 452192
rect 311866 452152 335360 452180
rect 335354 452140 335360 452152
rect 335412 452180 335418 452192
rect 336642 452180 336648 452192
rect 335412 452152 336648 452180
rect 335412 452140 335418 452152
rect 336642 452140 336648 452152
rect 336700 452140 336706 452192
rect 349706 452140 349712 452192
rect 349764 452180 349770 452192
rect 371234 452180 371240 452192
rect 349764 452152 371240 452180
rect 349764 452140 349770 452152
rect 371234 452140 371240 452152
rect 371292 452140 371298 452192
rect 378778 452140 378784 452192
rect 378836 452180 378842 452192
rect 385218 452180 385224 452192
rect 378836 452152 385224 452180
rect 378836 452140 378842 452152
rect 385218 452140 385224 452152
rect 385276 452140 385282 452192
rect 188246 452072 188252 452124
rect 188304 452112 188310 452124
rect 286502 452112 286508 452124
rect 188304 452084 286508 452112
rect 188304 452072 188310 452084
rect 286502 452072 286508 452084
rect 286560 452072 286566 452124
rect 291194 452072 291200 452124
rect 291252 452112 291258 452124
rect 297358 452112 297364 452124
rect 291252 452084 297364 452112
rect 291252 452072 291258 452084
rect 297358 452072 297364 452084
rect 297416 452072 297422 452124
rect 303982 452072 303988 452124
rect 304040 452112 304046 452124
rect 397178 452112 397184 452124
rect 304040 452084 397184 452112
rect 304040 452072 304046 452084
rect 397178 452072 397184 452084
rect 397236 452072 397242 452124
rect 191006 452004 191012 452056
rect 191064 452044 191070 452056
rect 290458 452044 290464 452056
rect 191064 452016 290464 452044
rect 191064 452004 191070 452016
rect 290458 452004 290464 452016
rect 290516 452004 290522 452056
rect 303890 452004 303896 452056
rect 303948 452044 303954 452056
rect 397086 452044 397092 452056
rect 303948 452016 397092 452044
rect 303948 452004 303954 452016
rect 397086 452004 397092 452016
rect 397144 452004 397150 452056
rect 189902 451936 189908 451988
rect 189960 451976 189966 451988
rect 295610 451976 295616 451988
rect 189960 451948 295616 451976
rect 189960 451936 189966 451948
rect 295610 451936 295616 451948
rect 295668 451976 295674 451988
rect 297634 451976 297640 451988
rect 295668 451948 297640 451976
rect 295668 451936 295674 451948
rect 297634 451936 297640 451948
rect 297692 451936 297698 451988
rect 297744 451948 303844 451976
rect 189994 451868 190000 451920
rect 190052 451908 190058 451920
rect 297744 451908 297772 451948
rect 190052 451880 297772 451908
rect 190052 451868 190058 451880
rect 297818 451868 297824 451920
rect 297876 451908 297882 451920
rect 303706 451908 303712 451920
rect 297876 451880 303712 451908
rect 297876 451868 297882 451880
rect 303706 451868 303712 451880
rect 303764 451868 303770 451920
rect 303816 451908 303844 451948
rect 304258 451936 304264 451988
rect 304316 451976 304322 451988
rect 396902 451976 396908 451988
rect 304316 451948 396908 451976
rect 304316 451936 304322 451948
rect 396902 451936 396908 451948
rect 396960 451936 396966 451988
rect 307754 451908 307760 451920
rect 303816 451880 307760 451908
rect 307754 451868 307760 451880
rect 307812 451908 307818 451920
rect 396994 451908 397000 451920
rect 307812 451880 397000 451908
rect 307812 451868 307818 451880
rect 396994 451868 397000 451880
rect 397052 451868 397058 451920
rect 191742 451800 191748 451852
rect 191800 451840 191806 451852
rect 314746 451840 314752 451852
rect 191800 451812 314752 451840
rect 191800 451800 191806 451812
rect 314746 451800 314752 451812
rect 314804 451800 314810 451852
rect 320818 451800 320824 451852
rect 320876 451840 320882 451852
rect 378778 451840 378784 451852
rect 320876 451812 378784 451840
rect 320876 451800 320882 451812
rect 378778 451800 378784 451812
rect 378836 451800 378842 451852
rect 380986 451800 380992 451852
rect 381044 451840 381050 451852
rect 381170 451840 381176 451852
rect 381044 451812 381176 451840
rect 381044 451800 381050 451812
rect 381170 451800 381176 451812
rect 381228 451800 381234 451852
rect 157794 451732 157800 451784
rect 157852 451772 157858 451784
rect 282362 451772 282368 451784
rect 157852 451744 282368 451772
rect 157852 451732 157858 451744
rect 282362 451732 282368 451744
rect 282420 451732 282426 451784
rect 297358 451732 297364 451784
rect 297416 451772 297422 451784
rect 394510 451772 394516 451784
rect 297416 451744 394516 451772
rect 297416 451732 297422 451744
rect 394510 451732 394516 451744
rect 394568 451732 394574 451784
rect 158622 451664 158628 451716
rect 158680 451704 158686 451716
rect 286410 451704 286416 451716
rect 158680 451676 286416 451704
rect 158680 451664 158686 451676
rect 286410 451664 286416 451676
rect 286468 451704 286474 451716
rect 413830 451704 413836 451716
rect 286468 451676 413836 451704
rect 286468 451664 286474 451676
rect 413830 451664 413836 451676
rect 413888 451664 413894 451716
rect 190914 451596 190920 451648
rect 190972 451636 190978 451648
rect 318794 451636 318800 451648
rect 190972 451608 318800 451636
rect 190972 451596 190978 451608
rect 318794 451596 318800 451608
rect 318852 451596 318858 451648
rect 336642 451596 336648 451648
rect 336700 451636 336706 451648
rect 388714 451636 388720 451648
rect 336700 451608 388720 451636
rect 336700 451596 336706 451608
rect 388714 451596 388720 451608
rect 388772 451596 388778 451648
rect 208302 451528 208308 451580
rect 208360 451568 208366 451580
rect 208578 451568 208584 451580
rect 208360 451540 208584 451568
rect 208360 451528 208366 451540
rect 208578 451528 208584 451540
rect 208636 451528 208642 451580
rect 253934 451528 253940 451580
rect 253992 451568 253998 451580
rect 254210 451568 254216 451580
rect 253992 451540 254216 451568
rect 253992 451528 253998 451540
rect 254210 451528 254216 451540
rect 254268 451528 254274 451580
rect 282362 451528 282368 451580
rect 282420 451568 282426 451580
rect 413738 451568 413744 451580
rect 282420 451540 413744 451568
rect 282420 451528 282426 451540
rect 413738 451528 413744 451540
rect 413796 451528 413802 451580
rect 158346 451460 158352 451512
rect 158404 451500 158410 451512
rect 282178 451500 282184 451512
rect 158404 451472 282184 451500
rect 158404 451460 158410 451472
rect 282178 451460 282184 451472
rect 282236 451460 282242 451512
rect 290826 451460 290832 451512
rect 290884 451500 290890 451512
rect 416498 451500 416504 451512
rect 290884 451472 416504 451500
rect 290884 451460 290890 451472
rect 416498 451460 416504 451472
rect 416556 451460 416562 451512
rect 156874 451392 156880 451444
rect 156932 451432 156938 451444
rect 299290 451432 299296 451444
rect 156932 451404 299296 451432
rect 156932 451392 156938 451404
rect 299290 451392 299296 451404
rect 299348 451392 299354 451444
rect 314746 451392 314752 451444
rect 314804 451432 314810 451444
rect 315482 451432 315488 451444
rect 314804 451404 315488 451432
rect 314804 451392 314810 451404
rect 315482 451392 315488 451404
rect 315540 451432 315546 451444
rect 320818 451432 320824 451444
rect 315540 451404 320824 451432
rect 315540 451392 315546 451404
rect 320818 451392 320824 451404
rect 320876 451392 320882 451444
rect 417418 451432 417424 451444
rect 325666 451404 417424 451432
rect 158438 451324 158444 451376
rect 158496 451364 158502 451376
rect 325418 451364 325424 451376
rect 158496 451336 325424 451364
rect 158496 451324 158502 451336
rect 325418 451324 325424 451336
rect 325476 451324 325482 451376
rect 187602 451256 187608 451308
rect 187660 451296 187666 451308
rect 196986 451296 196992 451308
rect 187660 451268 196992 451296
rect 187660 451256 187666 451268
rect 196986 451256 196992 451268
rect 197044 451256 197050 451308
rect 210510 451256 210516 451308
rect 210568 451296 210574 451308
rect 210568 451268 222332 451296
rect 210568 451256 210574 451268
rect 222304 451228 222332 451268
rect 222470 451256 222476 451308
rect 222528 451296 222534 451308
rect 222654 451296 222660 451308
rect 222528 451268 222660 451296
rect 222528 451256 222534 451268
rect 222654 451256 222660 451268
rect 222712 451256 222718 451308
rect 225690 451296 225696 451308
rect 223316 451268 225696 451296
rect 223316 451228 223344 451268
rect 225690 451256 225696 451268
rect 225748 451256 225754 451308
rect 278774 451256 278780 451308
rect 278832 451296 278838 451308
rect 296346 451296 296352 451308
rect 278832 451268 296352 451296
rect 278832 451256 278838 451268
rect 296346 451256 296352 451268
rect 296404 451256 296410 451308
rect 310514 451256 310520 451308
rect 310572 451296 310578 451308
rect 311802 451296 311808 451308
rect 310572 451268 311808 451296
rect 310572 451256 310578 451268
rect 311802 451256 311808 451268
rect 311860 451296 311866 451308
rect 325666 451296 325694 451404
rect 417418 451392 417424 451404
rect 417476 451392 417482 451444
rect 375190 451324 375196 451376
rect 375248 451364 375254 451376
rect 393038 451364 393044 451376
rect 375248 451336 393044 451364
rect 375248 451324 375254 451336
rect 393038 451324 393044 451336
rect 393096 451324 393102 451376
rect 311860 451268 325694 451296
rect 311860 451256 311866 451268
rect 373258 451256 373264 451308
rect 373316 451296 373322 451308
rect 419074 451296 419080 451308
rect 373316 451268 419080 451296
rect 373316 451256 373322 451268
rect 419074 451256 419080 451268
rect 419132 451256 419138 451308
rect 222304 451200 223344 451228
rect 166166 451052 166172 451104
rect 166224 451092 166230 451104
rect 350442 451092 350448 451104
rect 166224 451064 350448 451092
rect 166224 451052 166230 451064
rect 350442 451052 350448 451064
rect 350500 451052 350506 451104
rect 279418 450984 279424 451036
rect 279476 451024 279482 451036
rect 389818 451024 389824 451036
rect 279476 450996 389824 451024
rect 279476 450984 279482 450996
rect 389818 450984 389824 450996
rect 389876 450984 389882 451036
rect 280890 450916 280896 450968
rect 280948 450956 280954 450968
rect 409690 450956 409696 450968
rect 280948 450928 409696 450956
rect 280948 450916 280954 450928
rect 409690 450916 409696 450928
rect 409748 450916 409754 450968
rect 210418 450848 210424 450900
rect 210476 450888 210482 450900
rect 375098 450888 375104 450900
rect 210476 450860 375104 450888
rect 210476 450848 210482 450860
rect 375098 450848 375104 450860
rect 375156 450848 375162 450900
rect 191650 450780 191656 450832
rect 191708 450820 191714 450832
rect 281626 450820 281632 450832
rect 191708 450792 281632 450820
rect 191708 450780 191714 450792
rect 281626 450780 281632 450792
rect 281684 450780 281690 450832
rect 177942 450712 177948 450764
rect 178000 450752 178006 450764
rect 284570 450752 284576 450764
rect 178000 450724 284576 450752
rect 178000 450712 178006 450724
rect 284570 450712 284576 450724
rect 284628 450712 284634 450764
rect 298186 450712 298192 450764
rect 298244 450752 298250 450764
rect 298646 450752 298652 450764
rect 298244 450724 298652 450752
rect 298244 450712 298250 450724
rect 298646 450712 298652 450724
rect 298704 450712 298710 450764
rect 394602 450752 394608 450764
rect 302206 450724 394608 450752
rect 168190 450644 168196 450696
rect 168248 450684 168254 450696
rect 295242 450684 295248 450696
rect 168248 450656 295248 450684
rect 168248 450644 168254 450656
rect 295242 450644 295248 450656
rect 295300 450644 295306 450696
rect 298554 450644 298560 450696
rect 298612 450684 298618 450696
rect 302206 450684 302234 450724
rect 394602 450712 394608 450724
rect 394660 450712 394666 450764
rect 298612 450656 302234 450684
rect 298612 450644 298618 450656
rect 368842 450644 368848 450696
rect 368900 450684 368906 450696
rect 398558 450684 398564 450696
rect 368900 450656 398564 450684
rect 368900 450644 368906 450656
rect 398558 450644 398564 450656
rect 398616 450644 398622 450696
rect 3234 450576 3240 450628
rect 3292 450616 3298 450628
rect 210510 450616 210516 450628
rect 3292 450588 210516 450616
rect 3292 450576 3298 450588
rect 210510 450576 210516 450588
rect 210568 450576 210574 450628
rect 320634 450576 320640 450628
rect 320692 450616 320698 450628
rect 382182 450616 382188 450628
rect 320692 450588 382188 450616
rect 320692 450576 320698 450588
rect 382182 450576 382188 450588
rect 382240 450576 382246 450628
rect 17862 450508 17868 450560
rect 17920 450548 17926 450560
rect 278774 450548 278780 450560
rect 17920 450520 278780 450548
rect 17920 450508 17926 450520
rect 278774 450508 278780 450520
rect 278832 450508 278838 450560
rect 293770 450508 293776 450560
rect 293828 450548 293834 450560
rect 358722 450548 358728 450560
rect 293828 450520 358728 450548
rect 293828 450508 293834 450520
rect 358722 450508 358728 450520
rect 358780 450508 358786 450560
rect 365898 450508 365904 450560
rect 365956 450548 365962 450560
rect 401410 450548 401416 450560
rect 365956 450520 401416 450548
rect 365956 450508 365962 450520
rect 401410 450508 401416 450520
rect 401468 450508 401474 450560
rect 186130 450440 186136 450492
rect 186188 450480 186194 450492
rect 321738 450480 321744 450492
rect 186188 450452 321744 450480
rect 186188 450440 186194 450452
rect 321738 450440 321744 450452
rect 321796 450440 321802 450492
rect 365530 450440 365536 450492
rect 365588 450480 365594 450492
rect 409506 450480 409512 450492
rect 365588 450452 409512 450480
rect 365588 450440 365594 450452
rect 409506 450440 409512 450452
rect 409564 450440 409570 450492
rect 191558 450372 191564 450424
rect 191616 450412 191622 450424
rect 334986 450412 334992 450424
rect 191616 450384 334992 450412
rect 191616 450372 191622 450384
rect 334986 450372 334992 450384
rect 335044 450372 335050 450424
rect 336090 450372 336096 450424
rect 336148 450412 336154 450424
rect 403526 450412 403532 450424
rect 336148 450384 403532 450412
rect 336148 450372 336154 450384
rect 403526 450372 403532 450384
rect 403584 450372 403590 450424
rect 186038 450304 186044 450356
rect 186096 450344 186102 450356
rect 339770 450344 339776 450356
rect 186096 450316 339776 450344
rect 186096 450304 186102 450316
rect 339770 450304 339776 450316
rect 339828 450304 339834 450356
rect 346762 450304 346768 450356
rect 346820 450344 346826 450356
rect 395706 450344 395712 450356
rect 346820 450316 395712 450344
rect 346820 450304 346826 450316
rect 395706 450304 395712 450316
rect 395764 450304 395770 450356
rect 191834 450236 191840 450288
rect 191892 450276 191898 450288
rect 222102 450276 222108 450288
rect 191892 450248 222108 450276
rect 191892 450236 191898 450248
rect 222102 450236 222108 450248
rect 222160 450236 222166 450288
rect 222194 450236 222200 450288
rect 222252 450276 222258 450288
rect 222838 450276 222844 450288
rect 222252 450248 222844 450276
rect 222252 450236 222258 450248
rect 222838 450236 222844 450248
rect 222896 450236 222902 450288
rect 223574 450236 223580 450288
rect 223632 450276 223638 450288
rect 223942 450276 223948 450288
rect 223632 450248 223948 450276
rect 223632 450236 223638 450248
rect 223942 450236 223948 450248
rect 224000 450236 224006 450288
rect 244458 450236 244464 450288
rect 244516 450276 244522 450288
rect 245286 450276 245292 450288
rect 244516 450248 245292 450276
rect 244516 450236 244522 450248
rect 245286 450236 245292 450248
rect 245344 450236 245350 450288
rect 249794 450236 249800 450288
rect 249852 450276 249858 450288
rect 250070 450276 250076 450288
rect 249852 450248 250076 450276
rect 249852 450236 249858 450248
rect 250070 450236 250076 450248
rect 250128 450236 250134 450288
rect 252554 450236 252560 450288
rect 252612 450276 252618 450288
rect 252922 450276 252928 450288
rect 252612 450248 252928 450276
rect 252612 450236 252618 450248
rect 252922 450236 252928 450248
rect 252980 450236 252986 450288
rect 274726 450236 274732 450288
rect 274784 450276 274790 450288
rect 275094 450276 275100 450288
rect 274784 450248 275100 450276
rect 274784 450236 274790 450248
rect 275094 450236 275100 450248
rect 275152 450236 275158 450288
rect 302234 450236 302240 450288
rect 302292 450276 302298 450288
rect 302418 450276 302424 450288
rect 302292 450248 302424 450276
rect 302292 450236 302298 450248
rect 302418 450236 302424 450248
rect 302476 450236 302482 450288
rect 322934 450236 322940 450288
rect 322992 450276 322998 450288
rect 323302 450276 323308 450288
rect 322992 450248 323308 450276
rect 322992 450236 322998 450248
rect 323302 450236 323308 450248
rect 323360 450236 323366 450288
rect 362954 450236 362960 450288
rect 363012 450276 363018 450288
rect 363414 450276 363420 450288
rect 363012 450248 363420 450276
rect 363012 450236 363018 450248
rect 363414 450236 363420 450248
rect 363472 450236 363478 450288
rect 371418 450236 371424 450288
rect 371476 450276 371482 450288
rect 409414 450276 409420 450288
rect 371476 450248 409420 450276
rect 371476 450236 371482 450248
rect 409414 450236 409420 450248
rect 409472 450236 409478 450288
rect 177850 450168 177856 450220
rect 177908 450208 177914 450220
rect 351914 450208 351920 450220
rect 177908 450180 219434 450208
rect 177908 450168 177914 450180
rect 219406 450140 219434 450180
rect 222212 450180 351920 450208
rect 222212 450140 222240 450180
rect 351914 450168 351920 450180
rect 351972 450168 351978 450220
rect 362586 450168 362592 450220
rect 362644 450208 362650 450220
rect 412542 450208 412548 450220
rect 362644 450180 412548 450208
rect 362644 450168 362650 450180
rect 412542 450168 412548 450180
rect 412600 450168 412606 450220
rect 219406 450112 222240 450140
rect 222286 450100 222292 450152
rect 222344 450140 222350 450152
rect 227162 450140 227168 450152
rect 222344 450112 227168 450140
rect 222344 450100 222350 450112
rect 227162 450100 227168 450112
rect 227220 450100 227226 450152
rect 345290 450100 345296 450152
rect 345348 450140 345354 450152
rect 404262 450140 404268 450152
rect 345348 450112 404268 450140
rect 345348 450100 345354 450112
rect 404262 450100 404268 450112
rect 404320 450100 404326 450152
rect 165246 450032 165252 450084
rect 165304 450072 165310 450084
rect 290550 450072 290556 450084
rect 165304 450044 290556 450072
rect 165304 450032 165310 450044
rect 290550 450032 290556 450044
rect 290608 450032 290614 450084
rect 383470 450032 383476 450084
rect 383528 450072 383534 450084
rect 407022 450072 407028 450084
rect 383528 450044 407028 450072
rect 383528 450032 383534 450044
rect 407022 450032 407028 450044
rect 407080 450032 407086 450084
rect 3970 449964 3976 450016
rect 4028 450004 4034 450016
rect 226610 450004 226616 450016
rect 4028 449976 226616 450004
rect 4028 449964 4034 449976
rect 226610 449964 226616 449976
rect 226668 449964 226674 450016
rect 270494 449964 270500 450016
rect 270552 450004 270558 450016
rect 270770 450004 270776 450016
rect 270552 449976 270776 450004
rect 270552 449964 270558 449976
rect 270770 449964 270776 449976
rect 270828 449964 270834 450016
rect 325694 449964 325700 450016
rect 325752 450004 325758 450016
rect 325970 450004 325976 450016
rect 325752 449976 325976 450004
rect 325752 449964 325758 449976
rect 325970 449964 325976 449976
rect 326028 449964 326034 450016
rect 374270 449964 374276 450016
rect 374328 450004 374334 450016
rect 409598 450004 409604 450016
rect 374328 449976 409604 450004
rect 374328 449964 374334 449976
rect 409598 449964 409604 449976
rect 409656 449964 409662 450016
rect 19242 449896 19248 449948
rect 19300 449936 19306 449948
rect 278498 449936 278504 449948
rect 19300 449908 278504 449936
rect 19300 449896 19306 449908
rect 278498 449896 278504 449908
rect 278556 449896 278562 449948
rect 380802 449896 380808 449948
rect 380860 449936 380866 449948
rect 398466 449936 398472 449948
rect 380860 449908 398472 449936
rect 380860 449896 380866 449908
rect 398466 449896 398472 449908
rect 398524 449896 398530 449948
rect 190822 449828 190828 449880
rect 190880 449868 190886 449880
rect 193858 449868 193864 449880
rect 190880 449840 193864 449868
rect 190880 449828 190886 449840
rect 193858 449828 193864 449840
rect 193916 449828 193922 449880
rect 193950 449828 193956 449880
rect 194008 449868 194014 449880
rect 201218 449868 201224 449880
rect 194008 449840 201224 449868
rect 194008 449828 194014 449840
rect 201218 449828 201224 449840
rect 201276 449828 201282 449880
rect 198016 449772 202874 449800
rect 3694 449692 3700 449744
rect 3752 449732 3758 449744
rect 198016 449732 198044 449772
rect 3752 449704 198044 449732
rect 3752 449692 3758 449704
rect 200850 449692 200856 449744
rect 200908 449732 200914 449744
rect 202846 449732 202874 449772
rect 382274 449760 382280 449812
rect 382332 449800 382338 449812
rect 382332 449772 389174 449800
rect 382332 449760 382338 449772
rect 228082 449732 228088 449744
rect 200908 449704 201080 449732
rect 202846 449704 228088 449732
rect 200908 449692 200914 449704
rect 3878 449624 3884 449676
rect 3936 449664 3942 449676
rect 193122 449664 193128 449676
rect 3936 449636 193128 449664
rect 3936 449624 3942 449636
rect 193122 449624 193128 449636
rect 193180 449624 193186 449676
rect 193214 449624 193220 449676
rect 193272 449664 193278 449676
rect 195330 449664 195336 449676
rect 193272 449636 195336 449664
rect 193272 449624 193278 449636
rect 195330 449624 195336 449636
rect 195388 449624 195394 449676
rect 201052 449664 201080 449704
rect 228082 449692 228088 449704
rect 228140 449692 228146 449744
rect 382734 449692 382740 449744
rect 382792 449732 382798 449744
rect 386414 449732 386420 449744
rect 382792 449704 386420 449732
rect 382792 449692 382798 449704
rect 386414 449692 386420 449704
rect 386472 449692 386478 449744
rect 386506 449692 386512 449744
rect 386564 449732 386570 449744
rect 387610 449732 387616 449744
rect 386564 449704 387616 449732
rect 386564 449692 386570 449704
rect 387610 449692 387616 449704
rect 387668 449692 387674 449744
rect 387702 449692 387708 449744
rect 387760 449732 387766 449744
rect 388990 449732 388996 449744
rect 387760 449704 388996 449732
rect 387760 449692 387766 449704
rect 388990 449692 388996 449704
rect 389048 449692 389054 449744
rect 389146 449732 389174 449772
rect 413922 449732 413928 449744
rect 389146 449704 413928 449732
rect 413922 449692 413928 449704
rect 413980 449692 413986 449744
rect 201052 449636 202874 449664
rect 165338 449556 165344 449608
rect 165396 449596 165402 449608
rect 165396 449568 193214 449596
rect 165396 449556 165402 449568
rect 3510 449488 3516 449540
rect 3568 449528 3574 449540
rect 190822 449528 190828 449540
rect 3568 449500 190828 449528
rect 3568 449488 3574 449500
rect 190822 449488 190828 449500
rect 190880 449488 190886 449540
rect 193186 449528 193214 449568
rect 200850 449556 200856 449608
rect 200908 449556 200914 449608
rect 201218 449556 201224 449608
rect 201276 449556 201282 449608
rect 202846 449596 202874 449636
rect 379422 449624 379428 449676
rect 379480 449664 379486 449676
rect 416682 449664 416688 449676
rect 379480 449636 416688 449664
rect 379480 449624 379486 449636
rect 416682 449624 416688 449636
rect 416740 449624 416746 449676
rect 307202 449596 307208 449608
rect 202846 449568 307208 449596
rect 307202 449556 307208 449568
rect 307260 449556 307266 449608
rect 336734 449596 336740 449608
rect 316006 449568 336740 449596
rect 200868 449528 200896 449556
rect 193186 449500 200896 449528
rect 201236 449528 201264 449556
rect 316006 449528 316034 449568
rect 336734 449556 336740 449568
rect 336792 449556 336798 449608
rect 385218 449556 385224 449608
rect 385276 449556 385282 449608
rect 385678 449556 385684 449608
rect 385736 449596 385742 449608
rect 388070 449596 388076 449608
rect 385736 449568 388076 449596
rect 385736 449556 385742 449568
rect 388070 449556 388076 449568
rect 388128 449556 388134 449608
rect 399478 449596 399484 449608
rect 388180 449568 399484 449596
rect 201236 449500 316034 449528
rect 385236 449528 385264 449556
rect 388180 449528 388208 449568
rect 399478 449556 399484 449568
rect 399536 449556 399542 449608
rect 385236 449500 388208 449528
rect 388990 449488 388996 449540
rect 389048 449528 389054 449540
rect 411070 449528 411076 449540
rect 389048 449500 411076 449528
rect 389048 449488 389054 449500
rect 411070 449488 411076 449500
rect 411128 449488 411134 449540
rect 131758 444728 131764 444780
rect 131816 444768 131822 444780
rect 134334 444768 134340 444780
rect 131816 444740 134340 444768
rect 131816 444728 131822 444740
rect 134334 444728 134340 444740
rect 134392 444728 134398 444780
rect 151078 435344 151084 435396
rect 151136 435384 151142 435396
rect 158714 435384 158720 435396
rect 151136 435356 158720 435384
rect 151136 435344 151142 435356
rect 158714 435344 158720 435356
rect 158772 435344 158778 435396
rect 551922 435344 551928 435396
rect 551980 435384 551986 435396
rect 557534 435384 557540 435396
rect 551980 435356 557540 435384
rect 551980 435344 551986 435356
rect 557534 435344 557540 435356
rect 557592 435344 557598 435396
rect 19150 433984 19156 434036
rect 19208 434024 19214 434036
rect 131758 434024 131764 434036
rect 19208 433996 131764 434024
rect 19208 433984 19214 433996
rect 131758 433984 131764 433996
rect 131816 433984 131822 434036
rect 154574 433984 154580 434036
rect 154632 434024 154638 434036
rect 184198 434024 184204 434036
rect 154632 433996 184204 434024
rect 154632 433984 154638 433996
rect 184198 433984 184204 433996
rect 184256 433984 184262 434036
rect 558270 431876 558276 431928
rect 558328 431916 558334 431928
rect 580074 431916 580080 431928
rect 558328 431888 580080 431916
rect 558328 431876 558334 431888
rect 580074 431876 580080 431888
rect 580132 431876 580138 431928
rect 559558 419432 559564 419484
rect 559616 419472 559622 419484
rect 580074 419472 580080 419484
rect 559616 419444 580080 419472
rect 559616 419432 559622 419444
rect 580074 419432 580080 419444
rect 580132 419432 580138 419484
rect 563790 405628 563796 405680
rect 563848 405668 563854 405680
rect 580074 405668 580080 405680
rect 563848 405640 580080 405668
rect 563848 405628 563854 405640
rect 580074 405628 580080 405640
rect 580132 405628 580138 405680
rect 388898 384956 388904 385008
rect 388956 384996 388962 385008
rect 390370 384996 390376 385008
rect 388956 384968 390376 384996
rect 388956 384956 388962 384968
rect 390370 384956 390376 384968
rect 390428 384956 390434 385008
rect 17494 384276 17500 384328
rect 17552 384316 17558 384328
rect 18874 384316 18880 384328
rect 17552 384288 18880 384316
rect 17552 384276 17558 384288
rect 18874 384276 18880 384288
rect 18932 384276 18938 384328
rect 390278 382916 390284 382968
rect 390336 382956 390342 382968
rect 416774 382956 416780 382968
rect 390336 382928 416780 382956
rect 390336 382916 390342 382928
rect 416774 382916 416780 382928
rect 416832 382916 416838 382968
rect 17678 382236 17684 382288
rect 17736 382276 17742 382288
rect 18966 382276 18972 382288
rect 17736 382248 18972 382276
rect 17736 382236 17742 382248
rect 18966 382236 18972 382248
rect 19024 382236 19030 382288
rect 390186 381488 390192 381540
rect 390244 381528 390250 381540
rect 416866 381528 416872 381540
rect 390244 381500 416872 381528
rect 390244 381488 390250 381500
rect 416866 381488 416872 381500
rect 416924 381488 416930 381540
rect 390094 380128 390100 380180
rect 390152 380168 390158 380180
rect 416774 380168 416780 380180
rect 390152 380140 416780 380168
rect 390152 380128 390158 380140
rect 416774 380128 416780 380140
rect 416832 380128 416838 380180
rect 576118 379448 576124 379500
rect 576176 379488 576182 379500
rect 580074 379488 580080 379500
rect 576176 379460 580080 379488
rect 576176 379448 576182 379460
rect 580074 379448 580080 379460
rect 580132 379448 580138 379500
rect 388898 378768 388904 378820
rect 388956 378808 388962 378820
rect 416774 378808 416780 378820
rect 388956 378780 416780 378808
rect 388956 378768 388962 378780
rect 416774 378768 416780 378780
rect 416832 378768 416838 378820
rect 558178 353200 558184 353252
rect 558236 353240 558242 353252
rect 580074 353240 580080 353252
rect 558236 353212 580080 353240
rect 558236 353200 558242 353212
rect 580074 353200 580080 353212
rect 580132 353200 580138 353252
rect 399478 349868 399484 349920
rect 399536 349908 399542 349920
rect 418154 349908 418160 349920
rect 399536 349880 418160 349908
rect 399536 349868 399542 349880
rect 418154 349868 418160 349880
rect 418212 349868 418218 349920
rect 390370 349800 390376 349852
rect 390428 349840 390434 349852
rect 492582 349840 492588 349852
rect 390428 349812 492588 349840
rect 390428 349800 390434 349812
rect 492582 349800 492588 349812
rect 492640 349800 492646 349852
rect 103514 349596 103520 349648
rect 103572 349636 103578 349648
rect 162762 349636 162768 349648
rect 103572 349608 162768 349636
rect 103572 349596 103578 349608
rect 162762 349596 162768 349608
rect 162820 349596 162826 349648
rect 418154 349596 418160 349648
rect 418212 349636 418218 349648
rect 419442 349636 419448 349648
rect 418212 349608 419448 349636
rect 418212 349596 418218 349608
rect 419442 349596 419448 349608
rect 419500 349636 419506 349648
rect 452562 349636 452568 349648
rect 419500 349608 452568 349636
rect 419500 349596 419506 349608
rect 452562 349596 452568 349608
rect 452620 349596 452626 349648
rect 98546 349528 98552 349580
rect 98604 349568 98610 349580
rect 161290 349568 161296 349580
rect 98604 349540 161296 349568
rect 98604 349528 98610 349540
rect 161290 349528 161296 349540
rect 161348 349528 161354 349580
rect 408218 349528 408224 349580
rect 408276 349568 408282 349580
rect 478506 349568 478512 349580
rect 408276 349540 478512 349568
rect 408276 349528 408282 349540
rect 478506 349528 478512 349540
rect 478564 349528 478570 349580
rect 93486 349460 93492 349512
rect 93544 349500 93550 349512
rect 169662 349500 169668 349512
rect 93544 349472 169668 349500
rect 93544 349460 93550 349472
rect 169662 349460 169668 349472
rect 169720 349460 169726 349512
rect 400766 349460 400772 349512
rect 400824 349500 400830 349512
rect 483474 349500 483480 349512
rect 400824 349472 483480 349500
rect 400824 349460 400830 349472
rect 483474 349460 483480 349472
rect 483532 349460 483538 349512
rect 91002 349392 91008 349444
rect 91060 349432 91066 349444
rect 172330 349432 172336 349444
rect 91060 349404 172336 349432
rect 91060 349392 91066 349404
rect 172330 349392 172336 349404
rect 172388 349392 172394 349444
rect 398650 349392 398656 349444
rect 398708 349432 398714 349444
rect 485958 349432 485964 349444
rect 398708 349404 485964 349432
rect 398708 349392 398714 349404
rect 485958 349392 485964 349404
rect 486016 349392 486022 349444
rect 78030 349324 78036 349376
rect 78088 349364 78094 349376
rect 163406 349364 163412 349376
rect 78088 349336 163412 349364
rect 78088 349324 78094 349336
rect 163406 349324 163412 349336
rect 163464 349324 163470 349376
rect 395890 349324 395896 349376
rect 395948 349364 395954 349376
rect 488258 349364 488264 349376
rect 395948 349336 488264 349364
rect 395948 349324 395954 349336
rect 488258 349324 488264 349336
rect 488316 349324 488322 349376
rect 71774 349256 71780 349308
rect 71832 349296 71838 349308
rect 72234 349296 72240 349308
rect 71832 349268 72240 349296
rect 71832 349256 71838 349268
rect 72234 349256 72240 349268
rect 72292 349296 72298 349308
rect 190914 349296 190920 349308
rect 72292 349268 190920 349296
rect 72292 349256 72298 349268
rect 190914 349256 190920 349268
rect 190972 349256 190978 349308
rect 395798 349256 395804 349308
rect 395856 349296 395862 349308
rect 491018 349296 491024 349308
rect 395856 349268 491024 349296
rect 395856 349256 395862 349268
rect 491018 349256 491024 349268
rect 491076 349256 491082 349308
rect 67634 349188 67640 349240
rect 67692 349228 67698 349240
rect 68738 349228 68744 349240
rect 67692 349200 68744 349228
rect 67692 349188 67698 349200
rect 68738 349188 68744 349200
rect 68796 349228 68802 349240
rect 189994 349228 190000 349240
rect 68796 349200 190000 349228
rect 68796 349188 68802 349200
rect 189994 349188 190000 349200
rect 190052 349188 190058 349240
rect 416682 349188 416688 349240
rect 416740 349228 416746 349240
rect 520918 349228 520924 349240
rect 416740 349200 520924 349228
rect 416740 349188 416746 349200
rect 520918 349188 520924 349200
rect 520976 349188 520982 349240
rect 62850 349120 62856 349172
rect 62908 349160 62914 349172
rect 188246 349160 188252 349172
rect 62908 349132 188252 349160
rect 62908 349120 62914 349132
rect 188246 349120 188252 349132
rect 188304 349120 188310 349172
rect 393130 349120 393136 349172
rect 393188 349160 393194 349172
rect 508498 349160 508504 349172
rect 393188 349132 508504 349160
rect 393188 349120 393194 349132
rect 508498 349120 508504 349132
rect 508556 349120 508562 349172
rect 62022 349052 62028 349104
rect 62080 349092 62086 349104
rect 157794 349092 157800 349104
rect 62080 349064 157800 349092
rect 62080 349052 62086 349064
rect 157794 349052 157800 349064
rect 157852 349052 157858 349104
rect 388898 349052 388904 349104
rect 388956 349092 388962 349104
rect 419534 349092 419540 349104
rect 388956 349064 419540 349092
rect 388956 349052 388962 349064
rect 419534 349052 419540 349064
rect 419592 349052 419598 349104
rect 61102 348984 61108 349036
rect 61160 349024 61166 349036
rect 158530 349024 158536 349036
rect 61160 348996 158536 349024
rect 61160 348984 61166 348996
rect 158530 348984 158536 348996
rect 158588 348984 158594 349036
rect 414566 348984 414572 349036
rect 414624 349024 414630 349036
rect 418062 349024 418068 349036
rect 414624 348996 418068 349024
rect 414624 348984 414630 348996
rect 418062 348984 418068 348996
rect 418120 348984 418126 349036
rect 58526 348916 58532 348968
rect 58584 348956 58590 348968
rect 156874 348956 156880 348968
rect 58584 348928 156880 348956
rect 58584 348916 58590 348928
rect 156874 348916 156880 348928
rect 156932 348916 156938 348968
rect 56042 348848 56048 348900
rect 56100 348888 56106 348900
rect 156966 348888 156972 348900
rect 56100 348860 156972 348888
rect 56100 348848 56106 348860
rect 156966 348848 156972 348860
rect 157024 348848 157030 348900
rect 78490 348780 78496 348832
rect 78548 348820 78554 348832
rect 182726 348820 182732 348832
rect 78548 348792 182732 348820
rect 78548 348780 78554 348792
rect 182726 348780 182732 348792
rect 182784 348780 182790 348832
rect 419994 348780 420000 348832
rect 420052 348820 420058 348832
rect 500954 348820 500960 348832
rect 420052 348792 500960 348820
rect 420052 348780 420058 348792
rect 500954 348780 500960 348792
rect 501012 348780 501018 348832
rect 50798 348712 50804 348764
rect 50856 348752 50862 348764
rect 166902 348752 166908 348764
rect 50856 348724 166908 348752
rect 50856 348712 50862 348724
rect 166902 348712 166908 348724
rect 166960 348712 166966 348764
rect 418982 348712 418988 348764
rect 419040 348752 419046 348764
rect 505922 348752 505928 348764
rect 419040 348724 505928 348752
rect 419040 348712 419046 348724
rect 505922 348712 505928 348724
rect 505980 348712 505986 348764
rect 39574 348644 39580 348696
rect 39632 348684 39638 348696
rect 158622 348684 158628 348696
rect 39632 348656 158628 348684
rect 39632 348644 39638 348656
rect 158622 348644 158628 348656
rect 158680 348644 158686 348696
rect 411070 348644 411076 348696
rect 411128 348684 411134 348696
rect 418706 348684 418712 348696
rect 411128 348656 418712 348684
rect 411128 348644 411134 348656
rect 418706 348644 418712 348656
rect 418764 348644 418770 348696
rect 419074 348644 419080 348696
rect 419132 348684 419138 348696
rect 515858 348684 515864 348696
rect 419132 348656 515864 348684
rect 419132 348644 419138 348656
rect 515858 348644 515864 348656
rect 515916 348644 515922 348696
rect 38470 348576 38476 348628
rect 38528 348616 38534 348628
rect 158346 348616 158352 348628
rect 38528 348588 158352 348616
rect 38528 348576 38534 348588
rect 158346 348576 158352 348588
rect 158404 348576 158410 348628
rect 395614 348576 395620 348628
rect 395672 348616 395678 348628
rect 498470 348616 498476 348628
rect 395672 348588 498476 348616
rect 395672 348576 395678 348588
rect 498470 348576 498476 348588
rect 498528 348576 498534 348628
rect 71130 348508 71136 348560
rect 71188 348548 71194 348560
rect 190822 348548 190828 348560
rect 71188 348520 190828 348548
rect 71188 348508 71194 348520
rect 190822 348508 190828 348520
rect 190880 348508 190886 348560
rect 413922 348508 413928 348560
rect 413980 348548 413986 348560
rect 523310 348548 523316 348560
rect 413980 348520 523316 348548
rect 413980 348508 413986 348520
rect 523310 348508 523316 348520
rect 523368 348508 523374 348560
rect 65150 348440 65156 348492
rect 65208 348480 65214 348492
rect 189902 348480 189908 348492
rect 65208 348452 189908 348480
rect 65208 348440 65214 348452
rect 189902 348440 189908 348452
rect 189960 348440 189966 348492
rect 392946 348440 392952 348492
rect 393004 348480 393010 348492
rect 503438 348480 503444 348492
rect 393004 348452 503444 348480
rect 393004 348440 393010 348452
rect 503438 348440 503444 348452
rect 503496 348440 503502 348492
rect 53650 348372 53656 348424
rect 53708 348412 53714 348424
rect 190914 348412 190920 348424
rect 53708 348384 190920 348412
rect 53708 348372 53714 348384
rect 190914 348372 190920 348384
rect 190972 348372 190978 348424
rect 393038 348372 393044 348424
rect 393096 348412 393102 348424
rect 510982 348412 510988 348424
rect 393096 348384 510988 348412
rect 393096 348372 393102 348384
rect 510982 348372 510988 348384
rect 511040 348372 511046 348424
rect 86034 348304 86040 348356
rect 86092 348344 86098 348356
rect 177206 348344 177212 348356
rect 86092 348316 177212 348344
rect 86092 348304 86098 348316
rect 177206 348304 177212 348316
rect 177264 348304 177270 348356
rect 68370 348236 68376 348288
rect 68428 348276 68434 348288
rect 157886 348276 157892 348288
rect 68428 348248 157892 348276
rect 68428 348236 68434 348248
rect 157886 348236 157892 348248
rect 157944 348236 157950 348288
rect 73154 348168 73160 348220
rect 73212 348208 73218 348220
rect 74350 348208 74356 348220
rect 73212 348180 74356 348208
rect 73212 348168 73218 348180
rect 74350 348168 74356 348180
rect 74408 348208 74414 348220
rect 158438 348208 158444 348220
rect 74408 348180 158444 348208
rect 74408 348168 74414 348180
rect 158438 348168 158444 348180
rect 158496 348168 158502 348220
rect 418706 347896 418712 347948
rect 418764 347936 418770 347948
rect 455782 347936 455788 347948
rect 418764 347908 455788 347936
rect 418764 347896 418770 347908
rect 455782 347896 455788 347908
rect 455840 347896 455846 347948
rect 19150 347828 19156 347880
rect 19208 347868 19214 347880
rect 38470 347868 38476 347880
rect 19208 347840 38476 347868
rect 19208 347828 19214 347840
rect 38470 347828 38476 347840
rect 38528 347828 38534 347880
rect 419534 347828 419540 347880
rect 419592 347868 419598 347880
rect 458174 347868 458180 347880
rect 419592 347840 458180 347868
rect 419592 347828 419598 347840
rect 458174 347828 458180 347840
rect 458232 347828 458238 347880
rect 18690 347760 18696 347812
rect 18748 347800 18754 347812
rect 39574 347800 39580 347812
rect 18748 347772 39580 347800
rect 18748 347760 18754 347772
rect 39574 347760 39580 347772
rect 39632 347760 39638 347812
rect 418062 347760 418068 347812
rect 418120 347800 418126 347812
rect 456978 347800 456984 347812
rect 418120 347772 456984 347800
rect 418120 347760 418126 347772
rect 456978 347760 456984 347772
rect 457036 347800 457042 347812
rect 462222 347800 462228 347812
rect 457036 347772 462228 347800
rect 457036 347760 457042 347772
rect 462222 347760 462228 347772
rect 462280 347760 462286 347812
rect 42794 347692 42800 347744
rect 42852 347732 42858 347744
rect 62022 347732 62028 347744
rect 42852 347704 62028 347732
rect 42852 347692 42858 347704
rect 62022 347692 62028 347704
rect 62080 347692 62086 347744
rect 64782 347692 64788 347744
rect 64840 347732 64846 347744
rect 186958 347732 186964 347744
rect 64840 347704 186964 347732
rect 64840 347692 64846 347704
rect 186958 347692 186964 347704
rect 187016 347692 187022 347744
rect 417418 347692 417424 347744
rect 417476 347732 417482 347744
rect 417970 347732 417976 347744
rect 417476 347704 417976 347732
rect 417476 347692 417482 347704
rect 417970 347692 417976 347704
rect 418028 347692 418034 347744
rect 458174 347692 458180 347744
rect 458232 347732 458238 347744
rect 459462 347732 459468 347744
rect 458232 347704 459468 347732
rect 458232 347692 458238 347704
rect 459462 347692 459468 347704
rect 459520 347732 459526 347744
rect 478046 347732 478052 347744
rect 459520 347704 478052 347732
rect 459520 347692 459526 347704
rect 478046 347692 478052 347704
rect 478104 347692 478110 347744
rect 45922 347624 45928 347676
rect 45980 347664 45986 347676
rect 46566 347664 46572 347676
rect 45980 347636 46572 347664
rect 45980 347624 45986 347636
rect 46566 347624 46572 347636
rect 46624 347664 46630 347676
rect 65150 347664 65156 347676
rect 46624 347636 65156 347664
rect 46624 347624 46630 347636
rect 65150 347624 65156 347636
rect 65208 347624 65214 347676
rect 66254 347624 66260 347676
rect 66312 347664 66318 347676
rect 188890 347664 188896 347676
rect 66312 347636 188896 347664
rect 66312 347624 66318 347636
rect 188890 347624 188896 347636
rect 188948 347624 188954 347676
rect 394602 347624 394608 347676
rect 394660 347664 394666 347676
rect 458358 347664 458364 347676
rect 394660 347636 458364 347664
rect 394660 347624 394666 347636
rect 458358 347624 458364 347636
rect 458416 347624 458422 347676
rect 462222 347624 462228 347676
rect 462280 347664 462286 347676
rect 475654 347664 475660 347676
rect 462280 347636 475660 347664
rect 462280 347624 462286 347636
rect 475654 347624 475660 347636
rect 475712 347624 475718 347676
rect 477402 347624 477408 347676
rect 477460 347664 477466 347676
rect 479150 347664 479156 347676
rect 477460 347636 479156 347664
rect 477460 347624 477466 347636
rect 479150 347624 479156 347636
rect 479208 347624 479214 347676
rect 44174 347556 44180 347608
rect 44232 347596 44238 347608
rect 62850 347596 62856 347608
rect 44232 347568 62856 347596
rect 44232 347556 44238 347568
rect 62850 347556 62856 347568
rect 62908 347556 62914 347608
rect 67726 347556 67732 347608
rect 67784 347596 67790 347608
rect 187050 347596 187056 347608
rect 67784 347568 187056 347596
rect 67784 347556 67790 347568
rect 187050 347556 187056 347568
rect 187108 347556 187114 347608
rect 391382 347556 391388 347608
rect 391440 347596 391446 347608
rect 453574 347596 453580 347608
rect 391440 347568 453580 347596
rect 391440 347556 391446 347568
rect 453574 347556 453580 347568
rect 453632 347556 453638 347608
rect 455782 347556 455788 347608
rect 455840 347596 455846 347608
rect 474366 347596 474372 347608
rect 455840 347568 474372 347596
rect 455840 347556 455846 347568
rect 474366 347556 474372 347568
rect 474424 347556 474430 347608
rect 51074 347488 51080 347540
rect 51132 347528 51138 347540
rect 52362 347528 52368 347540
rect 51132 347500 52368 347528
rect 51132 347488 51138 347500
rect 52362 347488 52368 347500
rect 52420 347528 52426 347540
rect 71130 347528 71136 347540
rect 52420 347500 71136 347528
rect 52420 347488 52426 347500
rect 71130 347488 71136 347500
rect 71188 347488 71194 347540
rect 73246 347488 73252 347540
rect 73304 347528 73310 347540
rect 190822 347528 190828 347540
rect 73304 347500 190828 347528
rect 73304 347488 73310 347500
rect 190822 347488 190828 347500
rect 190880 347488 190886 347540
rect 391290 347488 391296 347540
rect 391348 347528 391354 347540
rect 450630 347528 450636 347540
rect 391348 347500 450636 347528
rect 391348 347488 391354 347500
rect 450630 347488 450636 347500
rect 450688 347488 450694 347540
rect 452562 347488 452568 347540
rect 452620 347528 452626 347540
rect 471238 347528 471244 347540
rect 452620 347500 471244 347528
rect 452620 347488 452626 347500
rect 471238 347488 471244 347500
rect 471296 347488 471302 347540
rect 53466 347460 53472 347472
rect 45526 347432 53472 347460
rect 16482 347216 16488 347268
rect 16540 347256 16546 347268
rect 45526 347256 45554 347432
rect 53466 347420 53472 347432
rect 53524 347460 53530 347472
rect 71774 347460 71780 347472
rect 53524 347432 71780 347460
rect 53524 347420 53530 347432
rect 71774 347420 71780 347432
rect 71832 347420 71838 347472
rect 76742 347420 76748 347472
rect 76800 347460 76806 347472
rect 190914 347460 190920 347472
rect 76800 347432 190920 347460
rect 76800 347420 76806 347432
rect 190914 347420 190920 347432
rect 190972 347420 190978 347472
rect 409690 347420 409696 347472
rect 409748 347460 409754 347472
rect 448238 347460 448244 347472
rect 409748 347432 448244 347460
rect 409748 347420 409754 347432
rect 448238 347420 448244 347432
rect 448296 347420 448302 347472
rect 50062 347352 50068 347404
rect 50120 347392 50126 347404
rect 67634 347392 67640 347404
rect 50120 347364 67640 347392
rect 50120 347352 50126 347364
rect 67634 347352 67640 347364
rect 67692 347352 67698 347404
rect 76098 347352 76104 347404
rect 76156 347392 76162 347404
rect 189810 347392 189816 347404
rect 76156 347364 189816 347392
rect 76156 347352 76162 347364
rect 189810 347352 189816 347364
rect 189868 347352 189874 347404
rect 416314 347352 416320 347404
rect 416372 347392 416378 347404
rect 418890 347392 418896 347404
rect 416372 347364 418896 347392
rect 416372 347352 416378 347364
rect 418890 347352 418896 347364
rect 418948 347352 418954 347404
rect 419350 347352 419356 347404
rect 419408 347392 419414 347404
rect 437014 347392 437020 347404
rect 419408 347364 437020 347392
rect 419408 347352 419414 347364
rect 437014 347352 437020 347364
rect 437072 347352 437078 347404
rect 73706 347284 73712 347336
rect 73764 347324 73770 347336
rect 186130 347324 186136 347336
rect 73764 347296 186136 347324
rect 73764 347284 73770 347296
rect 186130 347284 186136 347296
rect 186188 347284 186194 347336
rect 411806 347284 411812 347336
rect 411864 347324 411870 347336
rect 419718 347324 419724 347336
rect 411864 347296 419724 347324
rect 411864 347284 411870 347296
rect 419718 347284 419724 347296
rect 419776 347284 419782 347336
rect 436738 347284 436744 347336
rect 436796 347324 436802 347336
rect 443086 347324 443092 347336
rect 436796 347296 443092 347324
rect 436796 347284 436802 347296
rect 443086 347284 443092 347296
rect 443144 347324 443150 347336
rect 461486 347324 461492 347336
rect 443144 347296 461492 347324
rect 443144 347284 443150 347296
rect 461486 347284 461492 347296
rect 461544 347284 461550 347336
rect 16540 347228 45554 347256
rect 16540 347216 16546 347228
rect 56594 347216 56600 347268
rect 56652 347256 56658 347268
rect 73154 347256 73160 347268
rect 56652 347228 73160 347256
rect 56652 347216 56658 347228
rect 73154 347216 73160 347228
rect 73212 347216 73218 347268
rect 83642 347216 83648 347268
rect 83700 347256 83706 347268
rect 190822 347256 190828 347268
rect 83700 347228 190828 347256
rect 83700 347216 83706 347228
rect 190822 347216 190828 347228
rect 190880 347216 190886 347268
rect 413830 347216 413836 347268
rect 413888 347256 413894 347268
rect 419166 347256 419172 347268
rect 413888 347228 419172 347256
rect 413888 347216 413894 347228
rect 419166 347216 419172 347228
rect 419224 347216 419230 347268
rect 419258 347216 419264 347268
rect 419316 347256 419322 347268
rect 436094 347256 436100 347268
rect 419316 347228 436100 347256
rect 419316 347216 419322 347228
rect 436094 347216 436100 347228
rect 436152 347216 436158 347268
rect 452562 347216 452568 347268
rect 452620 347256 452626 347268
rect 469766 347256 469772 347268
rect 452620 347228 469772 347256
rect 452620 347216 452626 347228
rect 469766 347216 469772 347228
rect 469824 347216 469830 347268
rect 45370 347148 45376 347200
rect 45428 347188 45434 347200
rect 64782 347188 64788 347200
rect 45428 347160 64788 347188
rect 45428 347148 45434 347160
rect 19610 347080 19616 347132
rect 19668 347120 19674 347132
rect 37182 347120 37188 347132
rect 19668 347092 37188 347120
rect 19668 347080 19674 347092
rect 37182 347080 37188 347092
rect 37240 347080 37246 347132
rect 19886 347012 19892 347064
rect 19944 347052 19950 347064
rect 42794 347052 42800 347064
rect 19944 347024 42800 347052
rect 19944 347012 19950 347024
rect 42794 347012 42800 347024
rect 42852 347012 42858 347064
rect 19794 346944 19800 346996
rect 19852 346984 19858 346996
rect 44174 346984 44180 346996
rect 19852 346956 44180 346984
rect 19852 346944 19858 346956
rect 44174 346944 44180 346956
rect 44232 346944 44238 346996
rect 18966 346876 18972 346928
rect 19024 346916 19030 346928
rect 45526 346916 45554 347160
rect 64782 347148 64788 347160
rect 64840 347148 64846 347200
rect 81066 347148 81072 347200
rect 81124 347188 81130 347200
rect 179966 347188 179972 347200
rect 81124 347160 179972 347188
rect 81124 347148 81130 347160
rect 179966 347148 179972 347160
rect 180024 347148 180030 347200
rect 419074 347148 419080 347200
rect 419132 347188 419138 347200
rect 419132 347160 441614 347188
rect 419132 347148 419138 347160
rect 49602 347080 49608 347132
rect 49660 347120 49666 347132
rect 67726 347120 67732 347132
rect 49660 347092 67732 347120
rect 49660 347080 49666 347092
rect 67726 347080 67732 347092
rect 67784 347080 67790 347132
rect 100938 347080 100944 347132
rect 100996 347120 101002 347132
rect 190914 347120 190920 347132
rect 100996 347092 190920 347120
rect 100996 347080 101002 347092
rect 190914 347080 190920 347092
rect 190972 347080 190978 347132
rect 389910 347080 389916 347132
rect 389968 347120 389974 347132
rect 419626 347120 419632 347132
rect 389968 347092 419632 347120
rect 389968 347080 389974 347092
rect 419626 347080 419632 347092
rect 419684 347080 419690 347132
rect 419810 347080 419816 347132
rect 419868 347120 419874 347132
rect 440510 347120 440516 347132
rect 419868 347092 440516 347120
rect 419868 347080 419874 347092
rect 440510 347080 440516 347092
rect 440568 347080 440574 347132
rect 441586 347120 441614 347160
rect 456794 347148 456800 347200
rect 456852 347188 456858 347200
rect 458082 347188 458088 347200
rect 456852 347160 458088 347188
rect 456852 347148 456858 347160
rect 458082 347148 458088 347160
rect 458140 347188 458146 347200
rect 476942 347188 476948 347200
rect 458140 347160 476948 347188
rect 458140 347148 458146 347160
rect 476942 347148 476948 347160
rect 477000 347148 477006 347200
rect 444190 347120 444196 347132
rect 441586 347092 444196 347120
rect 444190 347080 444196 347092
rect 444248 347120 444254 347132
rect 462774 347120 462780 347132
rect 444248 347092 462780 347120
rect 444248 347080 444254 347092
rect 462774 347080 462780 347092
rect 462832 347080 462838 347132
rect 66254 347052 66260 347064
rect 19024 346888 45554 346916
rect 55186 347024 66260 347052
rect 19024 346876 19030 346888
rect 18598 346808 18604 346860
rect 18656 346848 18662 346860
rect 45922 346848 45928 346860
rect 18656 346820 45928 346848
rect 18656 346808 18662 346820
rect 45922 346808 45928 346820
rect 45980 346808 45986 346860
rect 16114 346740 16120 346792
rect 16172 346780 16178 346792
rect 47578 346780 47584 346792
rect 16172 346752 47584 346780
rect 16172 346740 16178 346752
rect 47578 346740 47584 346752
rect 47636 346780 47642 346792
rect 55186 346780 55214 347024
rect 66254 347012 66260 347024
rect 66312 347012 66318 347064
rect 75454 347012 75460 347064
rect 75512 347052 75518 347064
rect 162486 347052 162492 347064
rect 75512 347024 162492 347052
rect 75512 347012 75518 347024
rect 162486 347012 162492 347024
rect 162544 347012 162550 347064
rect 417970 347012 417976 347064
rect 418028 347052 418034 347064
rect 451366 347052 451372 347064
rect 418028 347024 451372 347052
rect 418028 347012 418034 347024
rect 451366 347012 451372 347024
rect 451424 347052 451430 347064
rect 452562 347052 452568 347064
rect 451424 347024 452568 347052
rect 451424 347012 451430 347024
rect 452562 347012 452568 347024
rect 452620 347012 452626 347064
rect 453022 347012 453028 347064
rect 453080 347052 453086 347064
rect 472066 347052 472072 347064
rect 453080 347024 472072 347052
rect 453080 347012 453086 347024
rect 472066 347012 472072 347024
rect 472124 347012 472130 347064
rect 60826 346944 60832 346996
rect 60884 346984 60890 346996
rect 78030 346984 78036 346996
rect 60884 346956 78036 346984
rect 60884 346944 60890 346956
rect 78030 346944 78036 346956
rect 78088 346944 78094 346996
rect 79134 346944 79140 346996
rect 79192 346984 79198 346996
rect 164142 346984 164148 346996
rect 79192 346956 164148 346984
rect 79192 346944 79198 346956
rect 164142 346944 164148 346956
rect 164200 346944 164206 346996
rect 391198 346944 391204 346996
rect 391256 346984 391262 346996
rect 456150 346984 456156 346996
rect 391256 346956 456156 346984
rect 391256 346944 391262 346956
rect 456150 346944 456156 346956
rect 456208 346944 456214 346996
rect 125962 346876 125968 346928
rect 126020 346916 126026 346928
rect 159818 346916 159824 346928
rect 126020 346888 159824 346916
rect 126020 346876 126026 346888
rect 159818 346876 159824 346888
rect 159876 346876 159882 346928
rect 416498 346876 416504 346928
rect 416556 346916 416562 346928
rect 419810 346916 419816 346928
rect 416556 346888 419816 346916
rect 416556 346876 416562 346888
rect 419810 346876 419816 346888
rect 419868 346876 419874 346928
rect 123386 346808 123392 346860
rect 123444 346848 123450 346860
rect 156690 346848 156696 346860
rect 123444 346820 156696 346848
rect 123444 346808 123450 346820
rect 156690 346808 156696 346820
rect 156748 346808 156754 346860
rect 419626 346808 419632 346860
rect 419684 346848 419690 346860
rect 456794 346848 456800 346860
rect 419684 346820 456800 346848
rect 419684 346808 419690 346820
rect 456794 346808 456800 346820
rect 456852 346808 456858 346860
rect 47636 346752 55214 346780
rect 47636 346740 47642 346752
rect 448514 346740 448520 346792
rect 448572 346780 448578 346792
rect 467374 346780 467380 346792
rect 448572 346752 467380 346780
rect 448572 346740 448578 346752
rect 467374 346740 467380 346752
rect 467432 346740 467438 346792
rect 18230 346672 18236 346724
rect 18288 346712 18294 346724
rect 18288 346684 50660 346712
rect 18288 346672 18294 346684
rect 16206 346604 16212 346656
rect 16264 346644 16270 346656
rect 48590 346644 48596 346656
rect 16264 346616 48596 346644
rect 16264 346604 16270 346616
rect 48590 346604 48596 346616
rect 48648 346644 48654 346656
rect 49602 346644 49608 346656
rect 48648 346616 49608 346644
rect 48648 346604 48654 346616
rect 49602 346604 49608 346616
rect 49660 346604 49666 346656
rect 16298 346536 16304 346588
rect 16356 346576 16362 346588
rect 50062 346576 50068 346588
rect 16356 346548 50068 346576
rect 16356 346536 16362 346548
rect 50062 346536 50068 346548
rect 50120 346536 50126 346588
rect 50632 346576 50660 346684
rect 55214 346672 55220 346724
rect 55272 346712 55278 346724
rect 73246 346712 73252 346724
rect 55272 346684 73252 346712
rect 55272 346672 55278 346684
rect 73246 346672 73252 346684
rect 73304 346672 73310 346724
rect 447134 346672 447140 346724
rect 447192 346712 447198 346724
rect 465718 346712 465724 346724
rect 447192 346684 465724 346712
rect 447192 346672 447198 346684
rect 465718 346672 465724 346684
rect 465776 346672 465782 346724
rect 59354 346604 59360 346656
rect 59412 346644 59418 346656
rect 76742 346644 76748 346656
rect 59412 346616 76748 346644
rect 59412 346604 59418 346616
rect 76742 346604 76748 346616
rect 76800 346604 76806 346656
rect 446398 346604 446404 346656
rect 446456 346644 446462 346656
rect 465166 346644 465172 346656
rect 446456 346616 465172 346644
rect 446456 346604 446462 346616
rect 465166 346604 465172 346616
rect 465224 346604 465230 346656
rect 51258 346576 51264 346588
rect 50632 346548 51264 346576
rect 51258 346536 51264 346548
rect 51316 346576 51322 346588
rect 69290 346576 69296 346588
rect 51316 346548 69296 346576
rect 51316 346536 51322 346548
rect 69290 346536 69296 346548
rect 69348 346536 69354 346588
rect 419166 346536 419172 346588
rect 419224 346576 419230 346588
rect 439590 346576 439596 346588
rect 419224 346548 439596 346576
rect 419224 346536 419230 346548
rect 439590 346536 439596 346548
rect 439648 346536 439654 346588
rect 445294 346536 445300 346588
rect 445352 346576 445358 346588
rect 463878 346576 463884 346588
rect 445352 346548 463884 346576
rect 445352 346536 445358 346548
rect 463878 346536 463884 346548
rect 463936 346536 463942 346588
rect 16390 346468 16396 346520
rect 16448 346508 16454 346520
rect 51074 346508 51080 346520
rect 16448 346480 51080 346508
rect 16448 346468 16454 346480
rect 51074 346468 51080 346480
rect 51132 346468 51138 346520
rect 61930 346468 61936 346520
rect 61988 346508 61994 346520
rect 79134 346508 79140 346520
rect 61988 346480 79140 346508
rect 61988 346468 61994 346480
rect 79134 346468 79140 346480
rect 79192 346468 79198 346520
rect 419718 346468 419724 346520
rect 419776 346508 419782 346520
rect 453022 346508 453028 346520
rect 419776 346480 453028 346508
rect 419776 346468 419782 346480
rect 453022 346468 453028 346480
rect 453080 346468 453086 346520
rect 455230 346468 455236 346520
rect 455288 346508 455294 346520
rect 473354 346508 473360 346520
rect 455288 346480 473360 346508
rect 455288 346468 455294 346480
rect 473354 346468 473360 346480
rect 473412 346468 473418 346520
rect 19702 346400 19708 346452
rect 19760 346440 19766 346452
rect 19760 346412 35894 346440
rect 19760 346400 19766 346412
rect 35866 346372 35894 346412
rect 418890 346400 418896 346452
rect 418948 346440 418954 346452
rect 438026 346440 438032 346452
rect 418948 346412 438032 346440
rect 418948 346400 418954 346412
rect 438026 346400 438032 346412
rect 438084 346400 438090 346452
rect 438854 346400 438860 346452
rect 438912 346440 438918 346452
rect 441614 346440 441620 346452
rect 438912 346412 441620 346440
rect 438912 346400 438918 346412
rect 441614 346400 441620 346412
rect 441672 346400 441678 346452
rect 449894 346400 449900 346452
rect 449952 346440 449958 346452
rect 468662 346440 468668 346452
rect 449952 346412 468668 346440
rect 449952 346400 449958 346412
rect 468662 346400 468668 346412
rect 468720 346400 468726 346452
rect 36170 346372 36176 346384
rect 35866 346344 36176 346372
rect 36170 346332 36176 346344
rect 36228 346372 36234 346384
rect 188982 346372 188988 346384
rect 36228 346344 188988 346372
rect 36228 346332 36234 346344
rect 188982 346332 188988 346344
rect 189040 346332 189046 346384
rect 394418 346332 394424 346384
rect 394476 346372 394482 346384
rect 525886 346372 525892 346384
rect 394476 346344 525892 346372
rect 394476 346332 394482 346344
rect 525886 346332 525892 346344
rect 525944 346332 525950 346384
rect 63678 346264 63684 346316
rect 63736 346304 63742 346316
rect 165338 346304 165344 346316
rect 63736 346276 165344 346304
rect 63736 346264 63742 346276
rect 165338 346264 165344 346276
rect 165396 346264 165402 346316
rect 392762 346264 392768 346316
rect 392820 346304 392826 346316
rect 518342 346304 518348 346316
rect 392820 346276 518348 346304
rect 392820 346264 392826 346276
rect 518342 346264 518348 346276
rect 518400 346264 518406 346316
rect 65978 346196 65984 346248
rect 66036 346236 66042 346248
rect 165062 346236 165068 346248
rect 66036 346208 165068 346236
rect 66036 346196 66042 346208
rect 165062 346196 165068 346208
rect 165120 346196 165126 346248
rect 392854 346196 392860 346248
rect 392912 346236 392918 346248
rect 513374 346236 513380 346248
rect 392912 346208 513380 346236
rect 392912 346196 392918 346208
rect 513374 346196 513380 346208
rect 513432 346196 513438 346248
rect 96062 346128 96068 346180
rect 96120 346168 96126 346180
rect 166166 346168 166172 346180
rect 96120 346140 166172 346168
rect 96120 346128 96126 346140
rect 166166 346128 166172 346140
rect 166224 346128 166230 346180
rect 394234 346128 394240 346180
rect 394292 346168 394298 346180
rect 465258 346168 465264 346180
rect 394292 346140 465264 346168
rect 394292 346128 394298 346140
rect 465258 346128 465264 346140
rect 465316 346128 465322 346180
rect 106090 346060 106096 346112
rect 106148 346100 106154 346112
rect 162394 346100 162400 346112
rect 106148 346072 162400 346100
rect 106148 346060 106154 346072
rect 162394 346060 162400 346072
rect 162452 346060 162458 346112
rect 413738 346060 413744 346112
rect 413796 346100 413802 346112
rect 419994 346100 420000 346112
rect 413796 346072 420000 346100
rect 413796 346060 413802 346072
rect 419994 346060 420000 346072
rect 420052 346060 420058 346112
rect 459554 346060 459560 346112
rect 459612 346100 459618 346112
rect 460566 346100 460572 346112
rect 459612 346072 460572 346100
rect 459612 346060 459618 346072
rect 460566 346060 460572 346072
rect 460624 346100 460630 346112
rect 477402 346100 477408 346112
rect 460624 346072 477408 346100
rect 460624 346060 460630 346072
rect 477402 346060 477408 346072
rect 477460 346060 477466 346112
rect 108666 345992 108672 346044
rect 108724 346032 108730 346044
rect 162302 346032 162308 346044
rect 108724 346004 162308 346032
rect 108724 345992 108730 346004
rect 162302 345992 162308 346004
rect 162360 345992 162366 346044
rect 394050 345992 394056 346044
rect 394108 346032 394114 346044
rect 460934 346032 460940 346044
rect 394108 346004 460940 346032
rect 394108 345992 394114 346004
rect 460934 345992 460940 346004
rect 460992 345992 460998 346044
rect 111058 345924 111064 345976
rect 111116 345964 111122 345976
rect 162578 345964 162584 345976
rect 111116 345936 162584 345964
rect 111116 345924 111122 345936
rect 162578 345924 162584 345936
rect 162636 345924 162642 345976
rect 396902 345924 396908 345976
rect 396960 345964 396966 345976
rect 414566 345964 414572 345976
rect 396960 345936 414572 345964
rect 396960 345924 396966 345936
rect 414566 345924 414572 345936
rect 414624 345964 414630 345976
rect 446398 345964 446404 345976
rect 414624 345936 446404 345964
rect 414624 345924 414630 345936
rect 446398 345924 446404 345936
rect 446456 345924 446462 345976
rect 115842 345856 115848 345908
rect 115900 345896 115906 345908
rect 165154 345896 165160 345908
rect 115900 345868 165160 345896
rect 115900 345856 115906 345868
rect 165154 345856 165160 345868
rect 165212 345856 165218 345908
rect 397178 345856 397184 345908
rect 397236 345896 397242 345908
rect 415854 345896 415860 345908
rect 397236 345868 415860 345896
rect 397236 345856 397242 345868
rect 415854 345856 415860 345868
rect 415912 345896 415918 345908
rect 448514 345896 448520 345908
rect 415912 345868 448520 345896
rect 415912 345856 415918 345868
rect 448514 345856 448520 345868
rect 448572 345856 448578 345908
rect 113450 345788 113456 345840
rect 113508 345828 113514 345840
rect 162670 345828 162676 345840
rect 113508 345800 162676 345828
rect 113508 345788 113514 345800
rect 162670 345788 162676 345800
rect 162728 345788 162734 345840
rect 394510 345788 394516 345840
rect 394568 345828 394574 345840
rect 415946 345828 415952 345840
rect 394568 345800 415952 345828
rect 394568 345788 394574 345800
rect 415946 345788 415952 345800
rect 416004 345788 416010 345840
rect 416682 345788 416688 345840
rect 416740 345828 416746 345840
rect 449894 345828 449900 345840
rect 416740 345800 449900 345828
rect 416740 345788 416746 345800
rect 449894 345788 449900 345800
rect 449952 345788 449958 345840
rect 118602 345720 118608 345772
rect 118660 345760 118666 345772
rect 164970 345760 164976 345772
rect 118660 345732 164976 345760
rect 118660 345720 118666 345732
rect 164970 345720 164976 345732
rect 165028 345720 165034 345772
rect 396810 345720 396816 345772
rect 396868 345760 396874 345772
rect 419902 345760 419908 345772
rect 396868 345732 419908 345760
rect 396868 345720 396874 345732
rect 419902 345720 419908 345732
rect 419960 345760 419966 345772
rect 455230 345760 455236 345772
rect 419960 345732 455236 345760
rect 419960 345720 419966 345732
rect 455230 345720 455236 345732
rect 455288 345720 455294 345772
rect 120994 345652 121000 345704
rect 121052 345692 121058 345704
rect 164878 345692 164884 345704
rect 121052 345664 164884 345692
rect 121052 345652 121058 345664
rect 164878 345652 164884 345664
rect 164936 345652 164942 345704
rect 396718 345652 396724 345704
rect 396776 345692 396782 345704
rect 414474 345692 414480 345704
rect 396776 345664 414480 345692
rect 396776 345652 396782 345664
rect 414474 345652 414480 345664
rect 414532 345692 414538 345704
rect 459554 345692 459560 345704
rect 414532 345664 459560 345692
rect 414532 345652 414538 345664
rect 459554 345652 459560 345664
rect 459612 345652 459618 345704
rect 397086 345584 397092 345636
rect 397144 345624 397150 345636
rect 416314 345624 416320 345636
rect 397144 345596 416320 345624
rect 397144 345584 397150 345596
rect 416314 345584 416320 345596
rect 416372 345624 416378 345636
rect 447134 345624 447140 345636
rect 416372 345596 447140 345624
rect 416372 345584 416378 345596
rect 447134 345584 447140 345596
rect 447192 345584 447198 345636
rect 415946 345516 415952 345568
rect 416004 345556 416010 345568
rect 445294 345556 445300 345568
rect 416004 345528 445300 345556
rect 416004 345516 416010 345528
rect 445294 345516 445300 345528
rect 445352 345516 445358 345568
rect 396994 345448 397000 345500
rect 397052 345488 397058 345500
rect 416682 345488 416688 345500
rect 397052 345460 416688 345488
rect 397052 345448 397058 345460
rect 416682 345448 416688 345460
rect 416740 345448 416746 345500
rect 419994 345448 420000 345500
rect 420052 345488 420058 345500
rect 436738 345488 436744 345500
rect 420052 345460 436744 345488
rect 420052 345448 420058 345460
rect 436738 345448 436744 345460
rect 436796 345448 436802 345500
rect 394326 345312 394332 345364
rect 394384 345352 394390 345364
rect 463510 345352 463516 345364
rect 394384 345324 463516 345352
rect 394384 345312 394390 345324
rect 463510 345312 463516 345324
rect 463568 345312 463574 345364
rect 19978 345040 19984 345092
rect 20036 345080 20042 345092
rect 41322 345080 41328 345092
rect 20036 345052 41328 345080
rect 20036 345040 20042 345052
rect 41322 345040 41328 345052
rect 41380 345040 41386 345092
rect 41340 344944 41368 345040
rect 42702 344972 42708 345024
rect 42760 345012 42766 345024
rect 168190 345012 168196 345024
rect 42760 344984 168196 345012
rect 42760 344972 42766 344984
rect 168190 344972 168196 344984
rect 168248 344972 168254 345024
rect 394142 344972 394148 345024
rect 394200 345012 394206 345024
rect 467926 345012 467932 345024
rect 394200 344984 467932 345012
rect 394200 344972 394206 344984
rect 467926 344972 467932 344984
rect 467984 344972 467990 345024
rect 165246 344944 165252 344956
rect 41340 344916 165252 344944
rect 165246 344904 165252 344916
rect 165304 344904 165310 344956
rect 69290 344836 69296 344888
rect 69348 344876 69354 344888
rect 168098 344876 168104 344888
rect 69348 344848 168104 344876
rect 69348 344836 69354 344848
rect 168098 344836 168104 344848
rect 168156 344836 168162 344888
rect 3418 344292 3424 344344
rect 3476 344332 3482 344344
rect 168006 344332 168012 344344
rect 3476 344304 168012 344332
rect 3476 344292 3482 344304
rect 168006 344292 168012 344304
rect 168064 344292 168070 344344
rect 418614 342932 418620 342984
rect 418672 342972 418678 342984
rect 418890 342972 418896 342984
rect 418672 342944 418896 342972
rect 418672 342932 418678 342944
rect 418890 342932 418896 342944
rect 418948 342932 418954 342984
rect 415854 340144 415860 340196
rect 415912 340184 415918 340196
rect 416498 340184 416504 340196
rect 415912 340156 416504 340184
rect 415912 340144 415918 340156
rect 416498 340144 416504 340156
rect 416556 340144 416562 340196
rect 551002 335452 551008 335504
rect 551060 335492 551066 335504
rect 557534 335492 557540 335504
rect 551060 335464 557540 335492
rect 551060 335452 551066 335464
rect 557534 335452 557540 335464
rect 557592 335452 557598 335504
rect 150986 335316 150992 335368
rect 151044 335356 151050 335368
rect 151044 335328 157380 335356
rect 151044 335316 151050 335328
rect 157352 335288 157380 335328
rect 158714 335288 158720 335300
rect 157352 335260 158720 335288
rect 158714 335248 158720 335260
rect 158772 335248 158778 335300
rect 18874 334908 18880 334960
rect 18932 334948 18938 334960
rect 55214 334948 55220 334960
rect 18932 334920 55220 334948
rect 18932 334908 18938 334920
rect 55214 334908 55220 334920
rect 55272 334908 55278 334960
rect 18322 334840 18328 334892
rect 18380 334880 18386 334892
rect 56594 334880 56600 334892
rect 18380 334852 56600 334880
rect 18380 334840 18386 334852
rect 56594 334840 56600 334852
rect 56652 334840 56658 334892
rect 18782 334772 18788 334824
rect 18840 334812 18846 334824
rect 57974 334812 57980 334824
rect 18840 334784 57980 334812
rect 18840 334772 18846 334784
rect 57974 334772 57980 334784
rect 58032 334772 58038 334824
rect 18506 334704 18512 334756
rect 18564 334744 18570 334756
rect 59354 334744 59360 334756
rect 18564 334716 59360 334744
rect 18564 334704 18570 334716
rect 59354 334704 59360 334716
rect 59412 334704 59418 334756
rect 19518 334636 19524 334688
rect 19576 334676 19582 334688
rect 60734 334676 60740 334688
rect 19576 334648 60740 334676
rect 19576 334636 19582 334648
rect 60734 334636 60740 334648
rect 60792 334636 60798 334688
rect 16022 334568 16028 334620
rect 16080 334608 16086 334620
rect 60826 334608 60832 334620
rect 16080 334580 60832 334608
rect 16080 334568 16086 334580
rect 60826 334568 60832 334580
rect 60884 334568 60890 334620
rect 563698 325592 563704 325644
rect 563756 325632 563762 325644
rect 579614 325632 579620 325644
rect 563756 325604 579620 325632
rect 563756 325592 563762 325604
rect 579614 325592 579620 325604
rect 579672 325592 579678 325644
rect 17034 259360 17040 259412
rect 17092 259400 17098 259412
rect 17310 259400 17316 259412
rect 17092 259372 17316 259400
rect 17092 259360 17098 259372
rect 17310 259360 17316 259372
rect 17368 259360 17374 259412
rect 392670 259360 392676 259412
rect 392728 259400 392734 259412
rect 417878 259400 417884 259412
rect 392728 259372 417884 259400
rect 392728 259360 392734 259372
rect 417878 259360 417884 259372
rect 417936 259360 417942 259412
rect 389910 258068 389916 258120
rect 389968 258108 389974 258120
rect 417142 258108 417148 258120
rect 389968 258080 417148 258108
rect 389968 258068 389974 258080
rect 417142 258068 417148 258080
rect 417200 258108 417206 258120
rect 418614 258108 418620 258120
rect 417200 258080 418620 258108
rect 417200 258068 417206 258080
rect 418614 258068 418620 258080
rect 418672 258068 418678 258120
rect 417694 253172 417700 253224
rect 417752 253212 417758 253224
rect 418614 253212 418620 253224
rect 417752 253184 418620 253212
rect 417752 253172 417758 253184
rect 418614 253172 418620 253184
rect 418672 253172 418678 253224
rect 388162 251812 388168 251864
rect 388220 251852 388226 251864
rect 406286 251852 406292 251864
rect 388220 251824 406292 251852
rect 388220 251812 388226 251824
rect 406286 251812 406292 251824
rect 406344 251812 406350 251864
rect 19334 249704 19340 249756
rect 19392 249744 19398 249756
rect 19610 249744 19616 249756
rect 19392 249716 19616 249744
rect 19392 249704 19398 249716
rect 19610 249704 19616 249716
rect 19668 249704 19674 249756
rect 111058 249704 111064 249756
rect 111116 249744 111122 249756
rect 174446 249744 174452 249756
rect 111116 249716 174452 249744
rect 111116 249704 111122 249716
rect 174446 249704 174452 249716
rect 174504 249704 174510 249756
rect 378226 249704 378232 249756
rect 378284 249744 378290 249756
rect 378778 249744 378784 249756
rect 378284 249716 378784 249744
rect 378284 249704 378290 249716
rect 378778 249704 378784 249716
rect 378836 249744 378842 249756
rect 389910 249744 389916 249756
rect 378836 249716 389916 249744
rect 378836 249704 378842 249716
rect 389910 249704 389916 249716
rect 389968 249704 389974 249756
rect 403526 249704 403532 249756
rect 403584 249744 403590 249756
rect 485958 249744 485964 249756
rect 403584 249716 485964 249744
rect 403584 249704 403590 249716
rect 485958 249704 485964 249716
rect 486016 249704 486022 249756
rect 108574 249636 108580 249688
rect 108632 249676 108638 249688
rect 174906 249676 174912 249688
rect 108632 249648 174912 249676
rect 108632 249636 108638 249648
rect 174906 249636 174912 249648
rect 174964 249636 174970 249688
rect 404170 249636 404176 249688
rect 404228 249676 404234 249688
rect 488258 249676 488264 249688
rect 404228 249648 488264 249676
rect 404228 249636 404234 249648
rect 488258 249636 488264 249648
rect 488316 249636 488322 249688
rect 19426 249568 19432 249620
rect 19484 249608 19490 249620
rect 19702 249608 19708 249620
rect 19484 249580 19708 249608
rect 19484 249568 19490 249580
rect 19702 249568 19708 249580
rect 19760 249568 19766 249620
rect 105998 249568 106004 249620
rect 106056 249608 106062 249620
rect 175182 249608 175188 249620
rect 106056 249580 175188 249608
rect 106056 249568 106062 249580
rect 175182 249568 175188 249580
rect 175240 249568 175246 249620
rect 404078 249568 404084 249620
rect 404136 249608 404142 249620
rect 491018 249608 491024 249620
rect 404136 249580 491024 249608
rect 404136 249568 404142 249580
rect 491018 249568 491024 249580
rect 491076 249568 491082 249620
rect 103514 249500 103520 249552
rect 103572 249540 103578 249552
rect 174814 249540 174820 249552
rect 103572 249512 174820 249540
rect 103572 249500 103578 249512
rect 174814 249500 174820 249512
rect 174872 249500 174878 249552
rect 401226 249500 401232 249552
rect 401284 249540 401290 249552
rect 495894 249540 495900 249552
rect 401284 249512 495900 249540
rect 401284 249500 401290 249512
rect 495894 249500 495900 249512
rect 495952 249500 495958 249552
rect 98546 249432 98552 249484
rect 98604 249472 98610 249484
rect 177850 249472 177856 249484
rect 98604 249444 177856 249472
rect 98604 249432 98610 249444
rect 177850 249432 177856 249444
rect 177908 249432 177914 249484
rect 401042 249432 401048 249484
rect 401100 249472 401106 249484
rect 498470 249472 498476 249484
rect 401100 249444 498476 249472
rect 401100 249432 401106 249444
rect 498470 249432 498476 249444
rect 498528 249432 498534 249484
rect 95878 249364 95884 249416
rect 95936 249404 95942 249416
rect 177482 249404 177488 249416
rect 95936 249376 177488 249404
rect 95936 249364 95942 249376
rect 177482 249364 177488 249376
rect 177540 249364 177546 249416
rect 308582 249364 308588 249416
rect 308640 249404 308646 249416
rect 311158 249404 311164 249416
rect 308640 249376 311164 249404
rect 308640 249364 308646 249376
rect 311158 249364 311164 249376
rect 311216 249364 311222 249416
rect 401134 249364 401140 249416
rect 401192 249404 401198 249416
rect 500954 249404 500960 249416
rect 401192 249376 500960 249404
rect 401192 249364 401198 249376
rect 500954 249364 500960 249376
rect 501012 249364 501018 249416
rect 93486 249296 93492 249348
rect 93544 249336 93550 249348
rect 177666 249336 177672 249348
rect 93544 249308 177672 249336
rect 93544 249296 93550 249308
rect 177666 249296 177672 249308
rect 177724 249296 177730 249348
rect 400950 249296 400956 249348
rect 401008 249336 401014 249348
rect 503530 249336 503536 249348
rect 401008 249308 503536 249336
rect 401008 249296 401014 249308
rect 503530 249296 503536 249308
rect 503588 249296 503594 249348
rect 58526 249228 58532 249280
rect 58584 249268 58590 249280
rect 172054 249268 172060 249280
rect 58584 249240 172060 249268
rect 58584 249228 58590 249240
rect 172054 249228 172060 249240
rect 172112 249228 172118 249280
rect 401502 249228 401508 249280
rect 401560 249268 401566 249280
rect 505922 249268 505928 249280
rect 401560 249240 505928 249268
rect 401560 249228 401566 249240
rect 505922 249228 505928 249240
rect 505980 249228 505986 249280
rect 56042 249160 56048 249212
rect 56100 249200 56106 249212
rect 172238 249200 172244 249212
rect 56100 249172 172244 249200
rect 56100 249160 56106 249172
rect 172238 249160 172244 249172
rect 172296 249160 172302 249212
rect 401318 249160 401324 249212
rect 401376 249200 401382 249212
rect 508498 249200 508504 249212
rect 401376 249172 508504 249200
rect 401376 249160 401382 249172
rect 508498 249160 508504 249172
rect 508556 249160 508562 249212
rect 53650 249092 53656 249144
rect 53708 249132 53714 249144
rect 172146 249132 172152 249144
rect 53708 249104 172152 249132
rect 53708 249092 53714 249104
rect 172146 249092 172152 249104
rect 172204 249092 172210 249144
rect 398190 249092 398196 249144
rect 398248 249132 398254 249144
rect 515858 249132 515864 249144
rect 398248 249104 515864 249132
rect 398248 249092 398254 249104
rect 515858 249092 515864 249104
rect 515916 249092 515922 249144
rect 15746 249024 15752 249076
rect 15804 249064 15810 249076
rect 18598 249064 18604 249076
rect 15804 249036 18604 249064
rect 15804 249024 15810 249036
rect 18598 249024 18604 249036
rect 18656 249064 18662 249076
rect 45922 249064 45928 249076
rect 18656 249036 45928 249064
rect 18656 249024 18662 249036
rect 45922 249024 45928 249036
rect 45980 249024 45986 249076
rect 50798 249024 50804 249076
rect 50856 249064 50862 249076
rect 177942 249064 177948 249076
rect 50856 249036 177948 249064
rect 50856 249024 50862 249036
rect 177942 249024 177948 249036
rect 178000 249024 178006 249076
rect 398282 249024 398288 249076
rect 398340 249064 398346 249076
rect 520918 249064 520924 249076
rect 398340 249036 520924 249064
rect 398340 249024 398346 249036
rect 520918 249024 520924 249036
rect 520976 249024 520982 249076
rect 113450 248956 113456 249008
rect 113508 248996 113514 249008
rect 174722 248996 174728 249008
rect 113508 248968 174728 248996
rect 113508 248956 113514 248968
rect 174722 248956 174728 248968
rect 174780 248956 174786 249008
rect 415302 248956 415308 249008
rect 415360 248996 415366 249008
rect 483474 248996 483480 249008
rect 415360 248968 483480 248996
rect 415360 248956 415366 248968
rect 483474 248956 483480 248968
rect 483532 248956 483538 249008
rect 115842 248888 115848 248940
rect 115900 248928 115906 248940
rect 174998 248928 175004 248940
rect 115900 248900 175004 248928
rect 115900 248888 115906 248900
rect 174998 248888 175004 248900
rect 175056 248888 175062 248940
rect 405366 248888 405372 248940
rect 405424 248928 405430 248940
rect 470962 248928 470968 248940
rect 405424 248900 470968 248928
rect 405424 248888 405430 248900
rect 470962 248888 470968 248900
rect 471020 248888 471026 248940
rect 120902 248820 120908 248872
rect 120960 248860 120966 248872
rect 174630 248860 174636 248872
rect 120960 248832 174636 248860
rect 120960 248820 120966 248832
rect 174630 248820 174636 248832
rect 174688 248820 174694 248872
rect 418798 248820 418804 248872
rect 418856 248860 418862 248872
rect 473630 248860 473636 248872
rect 418856 248832 473636 248860
rect 418856 248820 418862 248832
rect 473630 248820 473636 248832
rect 473688 248820 473694 248872
rect 19702 248452 19708 248464
rect 19444 248424 19708 248452
rect 16298 248344 16304 248396
rect 16356 248384 16362 248396
rect 19444 248384 19472 248424
rect 19702 248412 19708 248424
rect 19760 248452 19766 248464
rect 19760 248424 44220 248452
rect 19760 248412 19766 248424
rect 16356 248356 19472 248384
rect 44192 248384 44220 248424
rect 50154 248384 50160 248396
rect 44192 248356 50160 248384
rect 16356 248344 16362 248356
rect 50154 248344 50160 248356
rect 50212 248344 50218 248396
rect 61194 248344 61200 248396
rect 61252 248384 61258 248396
rect 171962 248384 171968 248396
rect 61252 248356 171968 248384
rect 61252 248344 61258 248356
rect 171962 248344 171968 248356
rect 172020 248344 172026 248396
rect 184198 248344 184204 248396
rect 184256 248384 184262 248396
rect 379606 248384 379612 248396
rect 184256 248356 379612 248384
rect 184256 248344 184262 248356
rect 379606 248344 379612 248356
rect 379664 248344 379670 248396
rect 382366 248344 382372 248396
rect 382424 248384 382430 248396
rect 382424 248356 384988 248384
rect 382424 248344 382430 248356
rect 19242 248276 19248 248328
rect 19300 248316 19306 248328
rect 36446 248316 36452 248328
rect 19300 248288 36452 248316
rect 19300 248276 19306 248288
rect 36446 248276 36452 248288
rect 36504 248276 36510 248328
rect 63586 248276 63592 248328
rect 63644 248316 63650 248328
rect 171870 248316 171876 248328
rect 63644 248288 171876 248316
rect 63644 248276 63650 248288
rect 171870 248276 171876 248288
rect 171928 248276 171934 248328
rect 18598 248208 18604 248260
rect 18656 248248 18662 248260
rect 19426 248248 19432 248260
rect 18656 248220 19432 248248
rect 18656 248208 18662 248220
rect 19426 248208 19432 248220
rect 19484 248248 19490 248260
rect 19484 248220 26234 248248
rect 19484 248208 19490 248220
rect 26206 248180 26234 248220
rect 29546 248208 29552 248260
rect 29604 248248 29610 248260
rect 38654 248248 38660 248260
rect 29604 248220 38660 248248
rect 29604 248208 29610 248220
rect 38654 248208 38660 248220
rect 38712 248208 38718 248260
rect 45922 248208 45928 248260
rect 45980 248248 45986 248260
rect 46658 248248 46664 248260
rect 45980 248220 46664 248248
rect 45980 248208 45986 248220
rect 46658 248208 46664 248220
rect 46716 248248 46722 248260
rect 64874 248248 64880 248260
rect 46716 248220 64880 248248
rect 46716 248208 46722 248220
rect 64874 248208 64880 248220
rect 64932 248208 64938 248260
rect 73798 248208 73804 248260
rect 73856 248248 73862 248260
rect 180518 248248 180524 248260
rect 73856 248220 180524 248248
rect 73856 248208 73862 248220
rect 180518 248208 180524 248220
rect 180576 248208 180582 248260
rect 384960 248248 384988 248356
rect 385126 248344 385132 248396
rect 385184 248384 385190 248396
rect 390646 248384 390652 248396
rect 385184 248356 390652 248384
rect 385184 248344 385190 248356
rect 390646 248344 390652 248356
rect 390704 248344 390710 248396
rect 402238 248276 402244 248328
rect 402296 248316 402302 248328
rect 455414 248316 455420 248328
rect 402296 248288 455420 248316
rect 402296 248276 402302 248288
rect 455414 248276 455420 248288
rect 455472 248276 455478 248328
rect 390554 248248 390560 248260
rect 384960 248220 390560 248248
rect 390554 248208 390560 248220
rect 390612 248208 390618 248260
rect 402330 248208 402336 248260
rect 402388 248248 402394 248260
rect 452654 248248 452660 248260
rect 402388 248220 452660 248248
rect 402388 248208 402394 248220
rect 452654 248208 452660 248220
rect 452712 248208 452718 248260
rect 35894 248180 35900 248192
rect 26206 248152 35900 248180
rect 35894 248140 35900 248152
rect 35952 248140 35958 248192
rect 44174 248140 44180 248192
rect 44232 248180 44238 248192
rect 62114 248180 62120 248192
rect 44232 248152 62120 248180
rect 44232 248140 44238 248152
rect 62114 248140 62120 248152
rect 62172 248140 62178 248192
rect 65978 248140 65984 248192
rect 66036 248180 66042 248192
rect 169478 248180 169484 248192
rect 66036 248152 169484 248180
rect 66036 248140 66042 248152
rect 169478 248140 169484 248152
rect 169536 248140 169542 248192
rect 383746 248140 383752 248192
rect 383804 248180 383810 248192
rect 390738 248180 390744 248192
rect 383804 248152 390744 248180
rect 383804 248140 383810 248152
rect 390738 248140 390744 248152
rect 390796 248140 390802 248192
rect 400858 248140 400864 248192
rect 400916 248180 400922 248192
rect 450354 248180 450360 248192
rect 400916 248152 450360 248180
rect 400916 248140 400922 248152
rect 450354 248140 450360 248152
rect 450412 248140 450418 248192
rect 19150 248072 19156 248124
rect 19208 248112 19214 248124
rect 37274 248112 37280 248124
rect 19208 248084 37280 248112
rect 19208 248072 19214 248084
rect 37274 248072 37280 248084
rect 37332 248072 37338 248124
rect 38102 248072 38108 248124
rect 38160 248112 38166 248124
rect 41414 248112 41420 248124
rect 38160 248084 41420 248112
rect 38160 248072 38166 248084
rect 41414 248072 41420 248084
rect 41472 248072 41478 248124
rect 59446 248072 59452 248124
rect 59504 248112 59510 248124
rect 77294 248112 77300 248124
rect 59504 248084 77300 248112
rect 59504 248072 59510 248084
rect 77294 248072 77300 248084
rect 77352 248072 77358 248124
rect 78490 248072 78496 248124
rect 78548 248112 78554 248124
rect 180610 248112 180616 248124
rect 78548 248084 180616 248112
rect 78548 248072 78554 248084
rect 180610 248072 180616 248084
rect 180668 248072 180674 248124
rect 380986 248072 380992 248124
rect 381044 248112 381050 248124
rect 389174 248112 389180 248124
rect 381044 248084 389180 248112
rect 381044 248072 381050 248084
rect 389174 248072 389180 248084
rect 389232 248072 389238 248124
rect 389818 248072 389824 248124
rect 389876 248112 389882 248124
rect 447134 248112 447140 248124
rect 389876 248084 447140 248112
rect 389876 248072 389882 248084
rect 447134 248072 447140 248084
rect 447192 248072 447198 248124
rect 450170 248072 450176 248124
rect 450228 248112 450234 248124
rect 451274 248112 451280 248124
rect 450228 248084 451280 248112
rect 450228 248072 450234 248084
rect 451274 248072 451280 248084
rect 451332 248112 451338 248124
rect 467834 248112 467840 248124
rect 451332 248084 467840 248112
rect 451332 248072 451338 248084
rect 467834 248072 467840 248084
rect 467892 248072 467898 248124
rect 19978 248004 19984 248056
rect 20036 248044 20042 248056
rect 40034 248044 40040 248056
rect 20036 248016 40040 248044
rect 20036 248004 20042 248016
rect 40034 248004 40040 248016
rect 40092 248004 40098 248056
rect 61378 248044 61384 248056
rect 43088 248016 61384 248044
rect 43088 247988 43116 248016
rect 61378 248004 61384 248016
rect 61436 248004 61442 248056
rect 68370 248004 68376 248056
rect 68428 248044 68434 248056
rect 169570 248044 169576 248056
rect 68428 248016 169576 248044
rect 68428 248004 68434 248016
rect 169570 248004 169576 248016
rect 169628 248004 169634 248056
rect 444466 248004 444472 248056
rect 444524 248044 444530 248056
rect 462314 248044 462320 248056
rect 444524 248016 462320 248044
rect 444524 248004 444530 248016
rect 462314 248004 462320 248016
rect 462372 248004 462378 248056
rect 19886 247936 19892 247988
rect 19944 247976 19950 247988
rect 43070 247976 43076 247988
rect 19944 247948 43076 247976
rect 19944 247936 19950 247948
rect 43070 247936 43076 247948
rect 43128 247936 43134 247988
rect 44266 247936 44272 247988
rect 44324 247976 44330 247988
rect 45278 247976 45284 247988
rect 44324 247948 45284 247976
rect 44324 247936 44330 247948
rect 45278 247936 45284 247948
rect 45336 247976 45342 247988
rect 63494 247976 63500 247988
rect 45336 247948 63500 247976
rect 45336 247936 45342 247948
rect 63494 247936 63500 247948
rect 63552 247936 63558 247988
rect 70946 247936 70952 247988
rect 71004 247976 71010 247988
rect 169386 247976 169392 247988
rect 71004 247948 169392 247976
rect 71004 247936 71010 247948
rect 169386 247936 169392 247948
rect 169444 247936 169450 247988
rect 443178 247936 443184 247988
rect 443236 247976 443242 247988
rect 444190 247976 444196 247988
rect 443236 247948 444196 247976
rect 443236 247936 443242 247948
rect 444190 247936 444196 247948
rect 444248 247976 444254 247988
rect 461118 247976 461124 247988
rect 444248 247948 461124 247976
rect 444248 247936 444254 247948
rect 461118 247936 461124 247948
rect 461176 247936 461182 247988
rect 19794 247868 19800 247920
rect 19852 247908 19858 247920
rect 44174 247908 44180 247920
rect 19852 247880 44180 247908
rect 19852 247868 19858 247880
rect 44174 247868 44180 247880
rect 44232 247868 44238 247920
rect 50154 247868 50160 247920
rect 50212 247908 50218 247920
rect 67634 247908 67640 247920
rect 50212 247880 67640 247908
rect 50212 247868 50218 247880
rect 67634 247868 67640 247880
rect 67692 247868 67698 247920
rect 83642 247868 83648 247920
rect 83700 247908 83706 247920
rect 180426 247908 180432 247920
rect 83700 247880 180432 247908
rect 83700 247868 83706 247880
rect 180426 247868 180432 247880
rect 180484 247868 180490 247920
rect 224218 247868 224224 247920
rect 224276 247908 224282 247920
rect 233326 247908 233332 247920
rect 224276 247880 233332 247908
rect 224276 247868 224282 247880
rect 233326 247868 233332 247880
rect 233384 247868 233390 247920
rect 447134 247868 447140 247920
rect 447192 247908 447198 247920
rect 465074 247908 465080 247920
rect 447192 247880 465080 247908
rect 447192 247868 447198 247880
rect 465074 247868 465080 247880
rect 465132 247868 465138 247920
rect 16114 247800 16120 247852
rect 16172 247840 16178 247852
rect 47578 247840 47584 247852
rect 16172 247812 47584 247840
rect 16172 247800 16178 247812
rect 47578 247800 47584 247812
rect 47636 247840 47642 247852
rect 66254 247840 66260 247852
rect 47636 247812 66260 247840
rect 47636 247800 47642 247812
rect 66254 247800 66260 247812
rect 66312 247800 66318 247852
rect 86034 247800 86040 247852
rect 86092 247840 86098 247852
rect 177758 247840 177764 247852
rect 86092 247812 177764 247840
rect 86092 247800 86098 247812
rect 177758 247800 177764 247812
rect 177816 247800 177822 247852
rect 220078 247800 220084 247852
rect 220136 247840 220142 247852
rect 229186 247840 229192 247852
rect 220136 247812 229192 247840
rect 220136 247800 220142 247812
rect 229186 247800 229192 247812
rect 229244 247800 229250 247852
rect 306466 247800 306472 247852
rect 306524 247840 306530 247852
rect 407114 247840 407120 247852
rect 306524 247812 407120 247840
rect 306524 247800 306530 247812
rect 407114 247800 407120 247812
rect 407172 247800 407178 247852
rect 451366 247800 451372 247852
rect 451424 247840 451430 247852
rect 452470 247840 452476 247852
rect 451424 247812 452476 247840
rect 451424 247800 451430 247812
rect 452470 247800 452476 247812
rect 452528 247840 452534 247852
rect 469214 247840 469220 247852
rect 452528 247812 469220 247840
rect 452528 247800 452534 247812
rect 469214 247800 469220 247812
rect 469272 247800 469278 247852
rect 16206 247732 16212 247784
rect 16264 247772 16270 247784
rect 48682 247772 48688 247784
rect 16264 247744 48688 247772
rect 16264 247732 16270 247744
rect 48682 247732 48688 247744
rect 48740 247772 48746 247784
rect 67726 247772 67732 247784
rect 48740 247744 67732 247772
rect 48740 247732 48746 247744
rect 67726 247732 67732 247744
rect 67784 247732 67790 247784
rect 88242 247732 88248 247784
rect 88300 247772 88306 247784
rect 177574 247772 177580 247784
rect 88300 247744 177580 247772
rect 88300 247732 88306 247744
rect 177574 247732 177580 247744
rect 177632 247732 177638 247784
rect 222838 247732 222844 247784
rect 222896 247772 222902 247784
rect 231946 247772 231952 247784
rect 222896 247744 231952 247772
rect 222896 247732 222902 247744
rect 231946 247732 231952 247744
rect 232004 247732 232010 247784
rect 307846 247732 307852 247784
rect 307904 247772 307910 247784
rect 409874 247772 409880 247784
rect 307904 247744 409880 247772
rect 307904 247732 307910 247744
rect 409874 247732 409880 247744
rect 409932 247732 409938 247784
rect 455874 247772 455880 247784
rect 451246 247744 455880 247772
rect 18506 247664 18512 247716
rect 18564 247704 18570 247716
rect 58066 247704 58072 247716
rect 18564 247676 58072 247704
rect 18564 247664 18570 247676
rect 58066 247664 58072 247676
rect 58124 247704 58130 247716
rect 75914 247704 75920 247716
rect 58124 247676 75920 247704
rect 58124 247664 58130 247676
rect 75914 247664 75920 247676
rect 75972 247664 75978 247716
rect 91002 247664 91008 247716
rect 91060 247704 91066 247716
rect 177298 247704 177304 247716
rect 91060 247676 177304 247704
rect 91060 247664 91066 247676
rect 177298 247664 177304 247676
rect 177356 247664 177362 247716
rect 218698 247664 218704 247716
rect 218756 247704 218762 247716
rect 227806 247704 227812 247716
rect 218756 247676 227812 247704
rect 218756 247664 218762 247676
rect 227806 247664 227812 247676
rect 227864 247664 227870 247716
rect 228358 247664 228364 247716
rect 228416 247704 228422 247716
rect 236086 247704 236092 247716
rect 228416 247676 236092 247704
rect 228416 247664 228422 247676
rect 236086 247664 236092 247676
rect 236144 247664 236150 247716
rect 309226 247664 309232 247716
rect 309284 247704 309290 247716
rect 414014 247704 414020 247716
rect 309284 247676 414020 247704
rect 309284 247664 309290 247676
rect 414014 247664 414020 247676
rect 414072 247664 414078 247716
rect 418522 247664 418528 247716
rect 418580 247704 418586 247716
rect 451246 247704 451274 247744
rect 455874 247732 455880 247744
rect 455932 247772 455938 247784
rect 473354 247772 473360 247784
rect 455932 247744 473360 247772
rect 455932 247732 455938 247744
rect 473354 247732 473360 247744
rect 473412 247732 473418 247784
rect 418580 247676 451274 247704
rect 418580 247664 418586 247676
rect 462222 247664 462228 247716
rect 462280 247704 462286 247716
rect 478874 247704 478880 247716
rect 462280 247676 478880 247704
rect 462280 247664 462286 247676
rect 478874 247664 478880 247676
rect 478932 247664 478938 247716
rect 15654 247596 15660 247648
rect 15712 247636 15718 247648
rect 18966 247636 18972 247648
rect 15712 247608 18972 247636
rect 15712 247596 15718 247608
rect 18966 247596 18972 247608
rect 19024 247636 19030 247648
rect 44266 247636 44272 247648
rect 19024 247608 44272 247636
rect 19024 247596 19030 247608
rect 44266 247596 44272 247608
rect 44324 247596 44330 247648
rect 63218 247596 63224 247648
rect 63276 247636 63282 247648
rect 74994 247636 75000 247648
rect 63276 247608 75000 247636
rect 63276 247596 63282 247608
rect 74994 247596 75000 247608
rect 75052 247596 75058 247648
rect 76098 247596 76104 247648
rect 76156 247636 76162 247648
rect 158254 247636 158260 247648
rect 76156 247608 158260 247636
rect 76156 247596 76162 247608
rect 158254 247596 158260 247608
rect 158312 247596 158318 247648
rect 449894 247596 449900 247648
rect 449952 247636 449958 247648
rect 466454 247636 466460 247648
rect 449952 247608 466460 247636
rect 449952 247596 449958 247608
rect 466454 247596 466460 247608
rect 466512 247596 466518 247648
rect 81066 247528 81072 247580
rect 81124 247568 81130 247580
rect 158070 247568 158076 247580
rect 81124 247540 158076 247568
rect 81124 247528 81130 247540
rect 158070 247528 158076 247540
rect 158128 247528 158134 247580
rect 448514 247528 448520 247580
rect 448572 247568 448578 247580
rect 465074 247568 465080 247580
rect 448572 247540 465080 247568
rect 448572 247528 448578 247540
rect 465074 247528 465080 247540
rect 465132 247528 465138 247580
rect 101214 247460 101220 247512
rect 101272 247500 101278 247512
rect 177390 247500 177396 247512
rect 101272 247472 177396 247500
rect 101272 247460 101278 247472
rect 177390 247460 177396 247472
rect 177448 247460 177454 247512
rect 452746 247460 452752 247512
rect 452804 247500 452810 247512
rect 470778 247500 470784 247512
rect 452804 247472 470784 247500
rect 452804 247460 452810 247472
rect 470778 247460 470784 247472
rect 470836 247460 470842 247512
rect 16022 247392 16028 247444
rect 16080 247432 16086 247444
rect 17034 247432 17040 247444
rect 16080 247404 17040 247432
rect 16080 247392 16086 247404
rect 17034 247392 17040 247404
rect 17092 247432 17098 247444
rect 59446 247432 59452 247444
rect 17092 247404 59452 247432
rect 17092 247392 17098 247404
rect 59446 247392 59452 247404
rect 59504 247392 59510 247444
rect 458266 247392 458272 247444
rect 458324 247432 458330 247444
rect 476114 247432 476120 247444
rect 458324 247404 476120 247432
rect 458324 247392 458330 247404
rect 476114 247392 476120 247404
rect 476172 247392 476178 247444
rect 52546 247324 52552 247376
rect 52604 247364 52610 247376
rect 69014 247364 69020 247376
rect 52604 247336 69020 247364
rect 52604 247324 52610 247336
rect 69014 247324 69020 247336
rect 69072 247324 69078 247376
rect 445754 247324 445760 247376
rect 445812 247364 445818 247376
rect 463694 247364 463700 247376
rect 445812 247336 463700 247364
rect 445812 247324 445818 247336
rect 463694 247324 463700 247336
rect 463752 247324 463758 247376
rect 52454 247256 52460 247308
rect 52512 247296 52518 247308
rect 70394 247296 70400 247308
rect 52512 247268 70400 247296
rect 52512 247256 52518 247268
rect 70394 247256 70400 247268
rect 70452 247256 70458 247308
rect 459554 247256 459560 247308
rect 459612 247296 459618 247308
rect 477494 247296 477500 247308
rect 459612 247268 477500 247296
rect 459612 247256 459618 247268
rect 477494 247256 477500 247268
rect 477552 247256 477558 247308
rect 53834 247188 53840 247240
rect 53892 247228 53898 247240
rect 71774 247228 71780 247240
rect 53892 247200 71780 247228
rect 53892 247188 53898 247200
rect 71774 247188 71780 247200
rect 71832 247188 71838 247240
rect 455414 247188 455420 247240
rect 455472 247228 455478 247240
rect 473354 247228 473360 247240
rect 455472 247200 473360 247228
rect 455472 247188 455478 247200
rect 473354 247188 473360 247200
rect 473412 247188 473418 247240
rect 18506 247120 18512 247172
rect 18564 247160 18570 247172
rect 19334 247160 19340 247172
rect 18564 247132 19340 247160
rect 18564 247120 18570 247132
rect 19334 247120 19340 247132
rect 19392 247120 19398 247172
rect 55122 247120 55128 247172
rect 55180 247160 55186 247172
rect 73154 247160 73160 247172
rect 55180 247132 73160 247160
rect 55180 247120 55186 247132
rect 73154 247120 73160 247132
rect 73212 247120 73218 247172
rect 454034 247120 454040 247172
rect 454092 247160 454098 247172
rect 471974 247160 471980 247172
rect 454092 247132 471980 247160
rect 454092 247120 454098 247132
rect 471974 247120 471980 247132
rect 472032 247120 472038 247172
rect 15930 247052 15936 247104
rect 15988 247092 15994 247104
rect 16206 247092 16212 247104
rect 15988 247064 16212 247092
rect 15988 247052 15994 247064
rect 16206 247052 16212 247064
rect 16264 247052 16270 247104
rect 19058 247052 19064 247104
rect 19116 247092 19122 247104
rect 19242 247092 19248 247104
rect 19116 247064 19248 247092
rect 19116 247052 19122 247064
rect 19242 247052 19248 247064
rect 19300 247052 19306 247104
rect 19426 247052 19432 247104
rect 19484 247092 19490 247104
rect 19978 247092 19984 247104
rect 19484 247064 19984 247092
rect 19484 247052 19490 247064
rect 19978 247052 19984 247064
rect 20036 247052 20042 247104
rect 56594 247052 56600 247104
rect 56652 247092 56658 247104
rect 73246 247092 73252 247104
rect 56652 247064 73252 247092
rect 56652 247052 56658 247064
rect 73246 247052 73252 247064
rect 73304 247052 73310 247104
rect 195238 247052 195244 247104
rect 195296 247092 195302 247104
rect 196066 247092 196072 247104
rect 195296 247064 196072 247092
rect 195296 247052 195302 247064
rect 196066 247052 196072 247064
rect 196124 247052 196130 247104
rect 199378 247052 199384 247104
rect 199436 247092 199442 247104
rect 200206 247092 200212 247104
rect 199436 247064 200212 247092
rect 199436 247052 199442 247064
rect 200206 247052 200212 247064
rect 200264 247052 200270 247104
rect 239398 247052 239404 247104
rect 239456 247092 239462 247104
rect 240226 247092 240232 247104
rect 239456 247064 240232 247092
rect 239456 247052 239462 247064
rect 240226 247052 240232 247064
rect 240284 247052 240290 247104
rect 271966 247052 271972 247104
rect 272024 247092 272030 247104
rect 273898 247092 273904 247104
rect 272024 247064 273904 247092
rect 272024 247052 272030 247064
rect 273898 247052 273904 247064
rect 273956 247052 273962 247104
rect 289906 247052 289912 247104
rect 289964 247092 289970 247104
rect 298738 247092 298744 247104
rect 289964 247064 298744 247092
rect 289964 247052 289970 247064
rect 298738 247052 298744 247064
rect 298796 247052 298802 247104
rect 299566 247052 299572 247104
rect 299624 247092 299630 247104
rect 302878 247092 302884 247104
rect 299624 247064 302884 247092
rect 299624 247052 299630 247064
rect 302878 247052 302884 247064
rect 302936 247052 302942 247104
rect 311986 247052 311992 247104
rect 312044 247092 312050 247104
rect 313918 247092 313924 247104
rect 312044 247064 313924 247092
rect 312044 247052 312050 247064
rect 313918 247052 313924 247064
rect 313976 247052 313982 247104
rect 325786 247052 325792 247104
rect 325844 247092 325850 247104
rect 329098 247092 329104 247104
rect 325844 247064 329104 247092
rect 325844 247052 325850 247064
rect 329098 247052 329104 247064
rect 329156 247052 329162 247104
rect 332686 247052 332692 247104
rect 332744 247092 332750 247104
rect 335998 247092 336004 247104
rect 332744 247064 336004 247092
rect 332744 247052 332750 247064
rect 335998 247052 336004 247064
rect 336056 247052 336062 247104
rect 398374 246984 398380 247036
rect 398432 247024 398438 247036
rect 525794 247024 525800 247036
rect 398432 246996 525800 247024
rect 398432 246984 398438 246996
rect 525794 246984 525800 246996
rect 525852 246984 525858 247036
rect 398558 246916 398564 246968
rect 398616 246956 398622 246968
rect 513374 246956 513380 246968
rect 398616 246928 513380 246956
rect 398616 246916 398622 246928
rect 513374 246916 513380 246928
rect 513432 246916 513438 246968
rect 401410 246848 401416 246900
rect 401468 246888 401474 246900
rect 510614 246888 510620 246900
rect 401468 246860 510620 246888
rect 401468 246848 401474 246860
rect 510614 246848 510620 246860
rect 510672 246848 510678 246900
rect 365806 246372 365812 246424
rect 365864 246412 365870 246424
rect 558178 246412 558184 246424
rect 365864 246384 558184 246412
rect 365864 246372 365870 246384
rect 558178 246372 558184 246384
rect 558236 246372 558242 246424
rect 372706 246304 372712 246356
rect 372764 246344 372770 246356
rect 576118 246344 576124 246356
rect 372764 246316 576124 246344
rect 372764 246304 372770 246316
rect 576118 246304 576124 246316
rect 576176 246304 576182 246356
rect 387058 245624 387064 245676
rect 387116 245664 387122 245676
rect 387886 245664 387892 245676
rect 387116 245636 387892 245664
rect 387116 245624 387122 245636
rect 387886 245624 387892 245636
rect 387944 245624 387950 245676
rect 398466 245556 398472 245608
rect 398524 245596 398530 245608
rect 523034 245596 523040 245608
rect 398524 245568 523040 245596
rect 398524 245556 398530 245568
rect 523034 245556 523040 245568
rect 523092 245556 523098 245608
rect 404262 245488 404268 245540
rect 404320 245528 404326 245540
rect 492674 245528 492680 245540
rect 404320 245500 492680 245528
rect 404320 245488 404326 245500
rect 492674 245488 492680 245500
rect 492732 245488 492738 245540
rect 403894 245420 403900 245472
rect 403952 245460 403958 245472
rect 480530 245460 480536 245472
rect 403952 245432 480536 245460
rect 403952 245420 403958 245432
rect 480530 245420 480536 245432
rect 480588 245420 480594 245472
rect 165614 244944 165620 244996
rect 165672 244984 165678 244996
rect 212626 244984 212632 244996
rect 165672 244956 212632 244984
rect 165672 244944 165678 244956
rect 212626 244944 212632 244956
rect 212684 244944 212690 244996
rect 7558 244876 7564 244928
rect 7616 244916 7622 244928
rect 191926 244916 191932 244928
rect 7616 244888 191932 244916
rect 7616 244876 7622 244888
rect 191926 244876 191932 244888
rect 191984 244876 191990 244928
rect 418614 243516 418620 243568
rect 418672 243556 418678 243568
rect 418982 243556 418988 243568
rect 418672 243528 418988 243556
rect 418672 243516 418678 243528
rect 418982 243516 418988 243528
rect 419040 243516 419046 243568
rect 186314 242156 186320 242208
rect 186372 242196 186378 242208
rect 220906 242196 220912 242208
rect 186372 242168 220912 242196
rect 186372 242156 186378 242168
rect 220906 242156 220912 242168
rect 220964 242156 220970 242208
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 167914 241448 167920 241460
rect 3568 241420 167920 241448
rect 3568 241408 3574 241420
rect 167914 241408 167920 241420
rect 167972 241408 167978 241460
rect 179414 240728 179420 240780
rect 179472 240768 179478 240780
rect 218054 240768 218060 240780
rect 179472 240740 218060 240768
rect 179472 240728 179478 240740
rect 218054 240728 218060 240740
rect 218112 240728 218118 240780
rect 387058 240728 387064 240780
rect 387116 240768 387122 240780
rect 557626 240768 557632 240780
rect 387116 240740 557632 240768
rect 387116 240728 387122 240740
rect 557626 240728 557632 240740
rect 557684 240768 557690 240780
rect 558822 240768 558828 240780
rect 557684 240740 558828 240768
rect 557684 240728 557690 240740
rect 558822 240728 558828 240740
rect 558880 240728 558886 240780
rect 419626 238688 419632 238740
rect 419684 238728 419690 238740
rect 458266 238728 458272 238740
rect 419684 238700 458272 238728
rect 419684 238688 419690 238700
rect 458266 238688 458272 238700
rect 458324 238688 458330 238740
rect 419810 238620 419816 238672
rect 419868 238660 419874 238672
rect 454034 238660 454040 238672
rect 419868 238632 454040 238660
rect 419868 238620 419874 238632
rect 454034 238620 454040 238632
rect 454092 238620 454098 238672
rect 368474 238076 368480 238128
rect 368532 238116 368538 238128
rect 562318 238116 562324 238128
rect 368532 238088 562324 238116
rect 368532 238076 368538 238088
rect 562318 238076 562324 238088
rect 562376 238076 562382 238128
rect 190178 238008 190184 238060
rect 190236 238048 190242 238060
rect 580534 238048 580540 238060
rect 190236 238020 580540 238048
rect 190236 238008 190242 238020
rect 580534 238008 580540 238020
rect 580592 238008 580598 238060
rect 415854 237396 415860 237448
rect 415912 237436 415918 237448
rect 419626 237436 419632 237448
rect 415912 237408 419632 237436
rect 415912 237396 415918 237408
rect 419626 237396 419632 237408
rect 419684 237396 419690 237448
rect 376754 236648 376760 236700
rect 376812 236688 376818 236700
rect 582374 236688 582380 236700
rect 376812 236660 582380 236688
rect 376812 236648 376818 236660
rect 582374 236648 582380 236660
rect 582432 236648 582438 236700
rect 17310 235900 17316 235952
rect 17368 235940 17374 235952
rect 150434 235940 150440 235952
rect 17368 235912 150440 235940
rect 17368 235900 17374 235912
rect 150434 235900 150440 235912
rect 150492 235900 150498 235952
rect 156690 235900 156696 235952
rect 156748 235940 156754 235952
rect 158622 235940 158628 235952
rect 156748 235912 158628 235940
rect 156748 235900 156754 235912
rect 158622 235900 158628 235912
rect 158680 235940 158686 235952
rect 378778 235940 378784 235952
rect 158680 235912 378784 235940
rect 158680 235900 158686 235912
rect 378778 235900 378784 235912
rect 378836 235900 378842 235952
rect 417694 235900 417700 235952
rect 417752 235940 417758 235952
rect 550818 235940 550824 235952
rect 417752 235912 550824 235940
rect 417752 235900 417758 235912
rect 550818 235900 550824 235912
rect 550876 235940 550882 235952
rect 557442 235940 557448 235952
rect 550876 235912 557448 235940
rect 550876 235900 550882 235912
rect 557442 235900 557448 235912
rect 557500 235900 557506 235952
rect 18322 235832 18328 235884
rect 18380 235872 18386 235884
rect 56594 235872 56600 235884
rect 18380 235844 56600 235872
rect 18380 235832 18386 235844
rect 56594 235832 56600 235844
rect 56652 235832 56658 235884
rect 418062 235832 418068 235884
rect 418120 235872 418126 235884
rect 458174 235872 458180 235884
rect 418120 235844 458180 235872
rect 418120 235832 418126 235844
rect 458174 235832 458180 235844
rect 458232 235832 458238 235884
rect 16298 235764 16304 235816
rect 16356 235804 16362 235816
rect 16482 235804 16488 235816
rect 16356 235776 16488 235804
rect 16356 235764 16362 235776
rect 16482 235764 16488 235776
rect 16540 235804 16546 235816
rect 53834 235804 53840 235816
rect 16540 235776 53840 235804
rect 16540 235764 16546 235776
rect 53834 235764 53840 235776
rect 53892 235764 53898 235816
rect 419902 235764 419908 235816
rect 419960 235804 419966 235816
rect 455414 235804 455420 235816
rect 419960 235776 455420 235804
rect 419960 235764 419966 235776
rect 455414 235764 455420 235776
rect 455472 235764 455478 235816
rect 16022 235696 16028 235748
rect 16080 235736 16086 235748
rect 16390 235736 16396 235748
rect 16080 235708 16396 235736
rect 16080 235696 16086 235708
rect 16390 235696 16396 235708
rect 16448 235736 16454 235748
rect 52454 235736 52460 235748
rect 16448 235708 52460 235736
rect 16448 235696 16454 235708
rect 52454 235696 52460 235708
rect 52512 235696 52518 235748
rect 416682 235696 416688 235748
rect 416740 235736 416746 235748
rect 451274 235736 451280 235748
rect 416740 235708 451280 235736
rect 416740 235696 416746 235708
rect 451274 235696 451280 235708
rect 451332 235696 451338 235748
rect 18874 235628 18880 235680
rect 18932 235668 18938 235680
rect 55214 235668 55220 235680
rect 18932 235640 55220 235668
rect 18932 235628 18938 235640
rect 55214 235628 55220 235640
rect 55272 235628 55278 235680
rect 416498 235628 416504 235680
rect 416556 235668 416562 235680
rect 449894 235668 449900 235680
rect 416556 235640 449900 235668
rect 416556 235628 416562 235640
rect 449894 235628 449900 235640
rect 449952 235628 449958 235680
rect 18230 235560 18236 235612
rect 18288 235600 18294 235612
rect 52546 235600 52552 235612
rect 18288 235572 52552 235600
rect 18288 235560 18294 235572
rect 52546 235560 52552 235572
rect 52604 235560 52610 235612
rect 419442 235560 419448 235612
rect 419500 235600 419506 235612
rect 452746 235600 452752 235612
rect 419500 235572 452752 235600
rect 419500 235560 419506 235572
rect 452746 235560 452752 235572
rect 452804 235560 452810 235612
rect 416314 235492 416320 235544
rect 416372 235532 416378 235544
rect 448514 235532 448520 235544
rect 416372 235504 448520 235532
rect 416372 235492 416378 235504
rect 448514 235492 448520 235504
rect 448572 235492 448578 235544
rect 419074 235424 419080 235476
rect 419132 235464 419138 235476
rect 444466 235464 444472 235476
rect 419132 235436 444472 235464
rect 419132 235424 419138 235436
rect 444466 235424 444472 235436
rect 444524 235424 444530 235476
rect 414566 235356 414572 235408
rect 414624 235396 414630 235408
rect 418982 235396 418988 235408
rect 414624 235368 418988 235396
rect 414624 235356 414630 235368
rect 418982 235356 418988 235368
rect 419040 235396 419046 235408
rect 447134 235396 447140 235408
rect 419040 235368 447140 235396
rect 419040 235356 419046 235368
rect 447134 235356 447140 235368
rect 447192 235356 447198 235408
rect 415946 235288 415952 235340
rect 416004 235328 416010 235340
rect 417142 235328 417148 235340
rect 416004 235300 417148 235328
rect 416004 235288 416010 235300
rect 417142 235288 417148 235300
rect 417200 235328 417206 235340
rect 445754 235328 445760 235340
rect 417200 235300 445760 235328
rect 417200 235288 417206 235300
rect 445754 235288 445760 235300
rect 445812 235288 445818 235340
rect 19518 235220 19524 235272
rect 19576 235260 19582 235272
rect 57974 235260 57980 235272
rect 19576 235232 57980 235260
rect 19576 235220 19582 235232
rect 57974 235220 57980 235232
rect 58032 235220 58038 235272
rect 311158 235220 311164 235272
rect 311216 235260 311222 235272
rect 340138 235260 340144 235272
rect 311216 235232 340144 235260
rect 311216 235220 311222 235232
rect 340138 235220 340144 235232
rect 340196 235220 340202 235272
rect 417970 235220 417976 235272
rect 418028 235260 418034 235272
rect 419534 235260 419540 235272
rect 418028 235232 419540 235260
rect 418028 235220 418034 235232
rect 419534 235220 419540 235232
rect 419592 235260 419598 235272
rect 452654 235260 452660 235272
rect 419592 235232 452660 235260
rect 419592 235220 419598 235232
rect 452654 235220 452660 235232
rect 452712 235220 452718 235272
rect 419718 235152 419724 235204
rect 419776 235192 419782 235204
rect 419994 235192 420000 235204
rect 419776 235164 420000 235192
rect 419776 235152 419782 235164
rect 419994 235152 420000 235164
rect 420052 235192 420058 235204
rect 444374 235192 444380 235204
rect 420052 235164 444380 235192
rect 420052 235152 420058 235164
rect 444374 235152 444380 235164
rect 444432 235152 444438 235204
rect 18230 235084 18236 235136
rect 18288 235124 18294 235136
rect 18690 235124 18696 235136
rect 18288 235096 18696 235124
rect 18288 235084 18294 235096
rect 18690 235084 18696 235096
rect 18748 235084 18754 235136
rect 418706 235084 418712 235136
rect 418764 235124 418770 235136
rect 419350 235124 419356 235136
rect 418764 235096 419356 235124
rect 418764 235084 418770 235096
rect 419350 235084 419356 235096
rect 419408 235124 419414 235136
rect 436094 235124 436100 235136
rect 419408 235096 436100 235124
rect 419408 235084 419414 235096
rect 436094 235084 436100 235096
rect 436152 235084 436158 235136
rect 418890 235016 418896 235068
rect 418948 235056 418954 235068
rect 419258 235056 419264 235068
rect 418948 235028 419264 235056
rect 418948 235016 418954 235028
rect 419258 235016 419264 235028
rect 419316 235056 419322 235068
rect 436186 235056 436192 235068
rect 419316 235028 436192 235056
rect 419316 235016 419322 235028
rect 436186 235016 436192 235028
rect 436244 235016 436250 235068
rect 18782 234948 18788 235000
rect 18840 234988 18846 235000
rect 19518 234988 19524 235000
rect 18840 234960 19524 234988
rect 18840 234948 18846 234960
rect 19518 234948 19524 234960
rect 19576 234948 19582 235000
rect 415670 234744 415676 234796
rect 415728 234784 415734 234796
rect 416498 234784 416504 234796
rect 415728 234756 416504 234784
rect 415728 234744 415734 234756
rect 416498 234744 416504 234756
rect 416556 234744 416562 234796
rect 415762 234676 415768 234728
rect 415820 234716 415826 234728
rect 416682 234716 416688 234728
rect 415820 234688 416688 234716
rect 415820 234676 415826 234688
rect 416682 234676 416688 234688
rect 416740 234676 416746 234728
rect 150434 234608 150440 234660
rect 150492 234648 150498 234660
rect 156690 234648 156696 234660
rect 150492 234620 156696 234648
rect 150492 234608 150498 234620
rect 156690 234608 156696 234620
rect 156748 234608 156754 234660
rect 416314 234608 416320 234660
rect 416372 234648 416378 234660
rect 416498 234648 416504 234660
rect 416372 234620 416504 234648
rect 416372 234608 416378 234620
rect 416498 234608 416504 234620
rect 416556 234608 416562 234660
rect 418430 234608 418436 234660
rect 418488 234648 418494 234660
rect 419074 234648 419080 234660
rect 418488 234620 419080 234648
rect 418488 234608 418494 234620
rect 419074 234608 419080 234620
rect 419132 234608 419138 234660
rect 556798 234540 556804 234592
rect 556856 234580 556862 234592
rect 557534 234580 557540 234592
rect 556856 234552 557540 234580
rect 556856 234540 556862 234552
rect 557534 234540 557540 234552
rect 557592 234540 557598 234592
rect 15838 233860 15844 233912
rect 15896 233900 15902 233912
rect 193214 233900 193220 233912
rect 15896 233872 193220 233900
rect 15896 233860 15902 233872
rect 193214 233860 193220 233872
rect 193272 233860 193278 233912
rect 197354 233860 197360 233912
rect 197412 233900 197418 233912
rect 224954 233900 224960 233912
rect 197412 233872 224960 233900
rect 197412 233860 197418 233872
rect 224954 233860 224960 233872
rect 225012 233860 225018 233912
rect 375374 233860 375380 233912
rect 375432 233900 375438 233912
rect 578878 233900 578884 233912
rect 375432 233872 578884 233900
rect 375432 233860 375438 233872
rect 578878 233860 578884 233872
rect 578936 233860 578942 233912
rect 577958 233180 577964 233232
rect 578016 233220 578022 233232
rect 579614 233220 579620 233232
rect 578016 233192 579620 233220
rect 578016 233180 578022 233192
rect 579614 233180 579620 233192
rect 579672 233180 579678 233232
rect 158714 230392 158720 230444
rect 158772 230432 158778 230444
rect 387058 230432 387064 230444
rect 158772 230404 387064 230432
rect 158772 230392 158778 230404
rect 387058 230392 387064 230404
rect 387116 230392 387122 230444
rect 172514 228352 172520 228404
rect 172572 228392 172578 228404
rect 215294 228392 215300 228404
rect 172572 228364 215300 228392
rect 172572 228352 172578 228364
rect 215294 228352 215300 228364
rect 215352 228352 215358 228404
rect 176654 226992 176660 227044
rect 176712 227032 176718 227044
rect 216674 227032 216680 227044
rect 176712 227004 216680 227032
rect 176712 226992 176718 227004
rect 216674 226992 216680 227004
rect 216732 226992 216738 227044
rect 303614 226992 303620 227044
rect 303672 227032 303678 227044
rect 398834 227032 398840 227044
rect 303672 227004 398840 227032
rect 303672 226992 303678 227004
rect 398834 226992 398840 227004
rect 398892 226992 398898 227044
rect 183554 225564 183560 225616
rect 183612 225604 183618 225616
rect 219434 225604 219440 225616
rect 183612 225576 219440 225604
rect 183612 225564 183618 225576
rect 219434 225564 219440 225576
rect 219492 225564 219498 225616
rect 340138 221076 340144 221128
rect 340196 221116 340202 221128
rect 345106 221116 345112 221128
rect 340196 221088 345112 221116
rect 340196 221076 340202 221088
rect 345106 221076 345112 221088
rect 345164 221076 345170 221128
rect 577866 219172 577872 219224
rect 577924 219212 577930 219224
rect 579982 219212 579988 219224
rect 577924 219184 579988 219212
rect 577924 219172 577930 219184
rect 579982 219172 579988 219184
rect 580040 219172 580046 219224
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 15102 215268 15108 215280
rect 3384 215240 15108 215268
rect 3384 215228 3390 215240
rect 15102 215228 15108 215240
rect 15160 215228 15166 215280
rect 345106 214548 345112 214600
rect 345164 214588 345170 214600
rect 359458 214588 359464 214600
rect 345164 214560 359464 214588
rect 345164 214548 345170 214560
rect 359458 214548 359464 214560
rect 359516 214548 359522 214600
rect 359458 207612 359464 207664
rect 359516 207652 359522 207664
rect 374638 207652 374644 207664
rect 359516 207624 374644 207652
rect 359516 207612 359522 207624
rect 374638 207612 374644 207624
rect 374696 207612 374702 207664
rect 273898 206252 273904 206304
rect 273956 206292 273962 206304
rect 317506 206292 317512 206304
rect 273956 206264 317512 206292
rect 273956 206252 273962 206264
rect 317506 206252 317512 206264
rect 317564 206252 317570 206304
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 15010 202824 15016 202836
rect 3108 202796 15016 202824
rect 3108 202784 3114 202796
rect 15010 202784 15016 202796
rect 15068 202784 15074 202836
rect 577774 193128 577780 193180
rect 577832 193168 577838 193180
rect 579614 193168 579620 193180
rect 577832 193140 579620 193168
rect 577832 193128 577838 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 14918 189020 14924 189032
rect 3568 188992 14924 189020
rect 3568 188980 3574 188992
rect 14918 188980 14924 188992
rect 14976 188980 14982 189032
rect 264974 180072 264980 180124
rect 265032 180112 265038 180124
rect 299474 180112 299480 180124
rect 265032 180084 299480 180112
rect 265032 180072 265038 180084
rect 299474 180072 299480 180084
rect 299532 180072 299538 180124
rect 302234 180072 302240 180124
rect 302292 180112 302298 180124
rect 396074 180112 396080 180124
rect 302292 180084 396080 180112
rect 302292 180072 302298 180084
rect 396074 180072 396080 180084
rect 396132 180072 396138 180124
rect 577682 179324 577688 179376
rect 577740 179364 577746 179376
rect 580074 179364 580080 179376
rect 577740 179336 580080 179364
rect 577740 179324 577746 179336
rect 580074 179324 580080 179336
rect 580132 179324 580138 179376
rect 260834 175924 260840 175976
rect 260892 175964 260898 175976
rect 287698 175964 287704 175976
rect 260892 175936 287704 175964
rect 260892 175924 260898 175936
rect 287698 175924 287704 175936
rect 287756 175924 287762 175976
rect 296714 175924 296720 175976
rect 296772 175964 296778 175976
rect 382274 175964 382280 175976
rect 296772 175936 382280 175964
rect 296772 175924 296778 175936
rect 382274 175924 382280 175936
rect 382332 175924 382338 175976
rect 374638 170280 374644 170332
rect 374696 170320 374702 170332
rect 377214 170320 377220 170332
rect 374696 170292 377220 170320
rect 374696 170280 374702 170292
rect 377214 170280 377220 170292
rect 377272 170280 377278 170332
rect 377214 167968 377220 168020
rect 377272 168008 377278 168020
rect 379514 168008 379520 168020
rect 377272 167980 379520 168008
rect 377272 167968 377278 167980
rect 379514 167968 379520 167980
rect 379572 167968 379578 168020
rect 379514 164840 379520 164892
rect 379572 164880 379578 164892
rect 400858 164880 400864 164892
rect 379572 164852 400864 164880
rect 379572 164840 379578 164852
rect 400858 164840 400864 164852
rect 400916 164840 400922 164892
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 14826 164200 14832 164212
rect 3292 164172 14832 164200
rect 3292 164160 3298 164172
rect 14826 164160 14832 164172
rect 14884 164160 14890 164212
rect 415210 158108 415216 158160
rect 415268 158148 415274 158160
rect 417694 158148 417700 158160
rect 415268 158120 417700 158148
rect 415268 158108 415274 158120
rect 417694 158108 417700 158120
rect 417752 158108 417758 158160
rect 400858 157972 400864 158024
rect 400916 158012 400922 158024
rect 410978 158012 410984 158024
rect 400916 157984 410984 158012
rect 400916 157972 400922 157984
rect 410978 157972 410984 157984
rect 411036 157972 411042 158024
rect 415854 149676 415860 149728
rect 415912 149716 415918 149728
rect 417694 149716 417700 149728
rect 415912 149688 417700 149716
rect 415912 149676 415918 149688
rect 417694 149676 417700 149688
rect 417752 149716 417758 149728
rect 458082 149716 458088 149728
rect 417752 149688 458088 149716
rect 417752 149676 417758 149688
rect 458082 149676 458088 149688
rect 458140 149676 458146 149728
rect 414750 149608 414756 149660
rect 414808 149648 414814 149660
rect 478506 149648 478512 149660
rect 414808 149620 478512 149648
rect 414808 149608 414814 149620
rect 478506 149608 478512 149620
rect 478564 149608 478570 149660
rect 415026 149540 415032 149592
rect 415084 149580 415090 149592
rect 480898 149580 480904 149592
rect 415084 149552 480904 149580
rect 415084 149540 415090 149552
rect 480898 149540 480904 149552
rect 480956 149540 480962 149592
rect 414842 149472 414848 149524
rect 414900 149512 414906 149524
rect 483474 149512 483480 149524
rect 414900 149484 483480 149512
rect 414900 149472 414906 149484
rect 483474 149472 483480 149484
rect 483532 149472 483538 149524
rect 412266 149404 412272 149456
rect 412324 149444 412330 149456
rect 485958 149444 485964 149456
rect 412324 149416 485964 149444
rect 412324 149404 412330 149416
rect 485958 149404 485964 149416
rect 486016 149404 486022 149456
rect 412450 149336 412456 149388
rect 412508 149376 412514 149388
rect 488258 149376 488264 149388
rect 412508 149348 488264 149376
rect 412508 149336 412514 149348
rect 488258 149336 488264 149348
rect 488316 149336 488322 149388
rect 412082 149268 412088 149320
rect 412140 149308 412146 149320
rect 491018 149308 491024 149320
rect 412140 149280 491024 149308
rect 412140 149268 412146 149280
rect 491018 149268 491024 149280
rect 491076 149268 491082 149320
rect 412174 149200 412180 149252
rect 412232 149240 412238 149252
rect 495894 149240 495900 149252
rect 412232 149212 495900 149240
rect 412232 149200 412238 149212
rect 495894 149200 495900 149212
rect 495952 149200 495958 149252
rect 412358 149132 412364 149184
rect 412416 149172 412422 149184
rect 503530 149172 503536 149184
rect 412416 149144 503536 149172
rect 412416 149132 412422 149144
rect 503530 149132 503536 149144
rect 503588 149132 503594 149184
rect 15102 149064 15108 149116
rect 15160 149104 15166 149116
rect 19610 149104 19616 149116
rect 15160 149076 19616 149104
rect 15160 149064 15166 149076
rect 19610 149064 19616 149076
rect 19668 149064 19674 149116
rect 409598 149064 409604 149116
rect 409656 149104 409662 149116
rect 518434 149104 518440 149116
rect 409656 149076 518440 149104
rect 409656 149064 409662 149076
rect 518434 149064 518440 149076
rect 518492 149064 518498 149116
rect 98546 148996 98552 149048
rect 98604 149036 98610 149048
rect 183462 149036 183468 149048
rect 98604 149008 183468 149036
rect 98604 148996 98610 149008
rect 183462 148996 183468 149008
rect 183520 148996 183526 149048
rect 403710 148996 403716 149048
rect 403768 149036 403774 149048
rect 468294 149036 468300 149048
rect 403768 149008 468300 149036
rect 403768 148996 403774 149008
rect 468294 148996 468300 149008
rect 468352 148996 468358 149048
rect 93486 148928 93492 148980
rect 93544 148968 93550 148980
rect 185946 148968 185952 148980
rect 93544 148940 185952 148968
rect 93544 148928 93550 148940
rect 185946 148928 185952 148940
rect 186004 148928 186010 148980
rect 403802 148928 403808 148980
rect 403860 148968 403866 148980
rect 470962 148968 470968 148980
rect 403860 148940 470968 148968
rect 403860 148928 403866 148940
rect 470962 148928 470968 148940
rect 471020 148928 471026 148980
rect 86034 148860 86040 148912
rect 86092 148900 86098 148912
rect 185670 148900 185676 148912
rect 86092 148872 185676 148900
rect 86092 148860 86098 148872
rect 185670 148860 185676 148872
rect 185728 148860 185734 148912
rect 411990 148860 411996 148912
rect 412048 148900 412054 148912
rect 505922 148900 505928 148912
rect 412048 148872 505928 148900
rect 412048 148860 412054 148872
rect 505922 148860 505928 148872
rect 505980 148860 505986 148912
rect 83550 148792 83556 148844
rect 83608 148832 83614 148844
rect 188706 148832 188712 148844
rect 83608 148804 188712 148832
rect 83608 148792 83614 148804
rect 188706 148792 188712 148804
rect 188764 148792 188770 148844
rect 412542 148792 412548 148844
rect 412600 148832 412606 148844
rect 508498 148832 508504 148844
rect 412600 148804 508504 148832
rect 412600 148792 412606 148804
rect 508498 148792 508504 148804
rect 508556 148792 508562 148844
rect 76098 148724 76104 148776
rect 76156 148764 76162 148776
rect 188614 148764 188620 148776
rect 76156 148736 188620 148764
rect 76156 148724 76162 148736
rect 188614 148724 188620 148736
rect 188672 148724 188678 148776
rect 409506 148724 409512 148776
rect 409564 148764 409570 148776
rect 510982 148764 510988 148776
rect 409564 148736 510988 148764
rect 409564 148724 409570 148736
rect 510982 148724 510988 148736
rect 511040 148724 511046 148776
rect 19610 148656 19616 148708
rect 19668 148696 19674 148708
rect 60642 148696 60648 148708
rect 19668 148668 60648 148696
rect 19668 148656 19674 148668
rect 60642 148656 60648 148668
rect 60700 148656 60706 148708
rect 73614 148656 73620 148708
rect 73672 148696 73678 148708
rect 188522 148696 188528 148708
rect 73672 148668 188528 148696
rect 73672 148656 73678 148668
rect 188522 148656 188528 148668
rect 188580 148656 188586 148708
rect 409230 148656 409236 148708
rect 409288 148696 409294 148708
rect 513374 148696 513380 148708
rect 409288 148668 513380 148696
rect 409288 148656 409294 148668
rect 513374 148656 513380 148668
rect 513432 148656 513438 148708
rect 58526 148588 58532 148640
rect 58584 148628 58590 148640
rect 180242 148628 180248 148640
rect 58584 148600 180248 148628
rect 58584 148588 58590 148600
rect 180242 148588 180248 148600
rect 180300 148588 180306 148640
rect 409414 148588 409420 148640
rect 409472 148628 409478 148640
rect 515858 148628 515864 148640
rect 409472 148600 515864 148628
rect 409472 148588 409478 148600
rect 515858 148588 515864 148600
rect 515916 148588 515922 148640
rect 56042 148520 56048 148572
rect 56100 148560 56106 148572
rect 180334 148560 180340 148572
rect 56100 148532 180340 148560
rect 56100 148520 56106 148532
rect 180334 148520 180340 148532
rect 180392 148520 180398 148572
rect 409322 148520 409328 148572
rect 409380 148560 409386 148572
rect 520918 148560 520924 148572
rect 409380 148532 520924 148560
rect 409380 148520 409386 148532
rect 520918 148520 520924 148532
rect 520976 148520 520982 148572
rect 53650 148452 53656 148504
rect 53708 148492 53714 148504
rect 183278 148492 183284 148504
rect 53708 148464 183284 148492
rect 53708 148452 53714 148464
rect 183278 148452 183284 148464
rect 183336 148452 183342 148504
rect 406930 148452 406936 148504
rect 406988 148492 406994 148504
rect 523310 148492 523316 148504
rect 406988 148464 523316 148492
rect 406988 148452 406994 148464
rect 523310 148452 523316 148464
rect 523368 148452 523374 148504
rect 19702 148384 19708 148436
rect 19760 148424 19766 148436
rect 19978 148424 19984 148436
rect 19760 148396 19984 148424
rect 19760 148384 19766 148396
rect 19978 148384 19984 148396
rect 20036 148384 20042 148436
rect 50798 148384 50804 148436
rect 50856 148424 50862 148436
rect 185854 148424 185860 148436
rect 50856 148396 185860 148424
rect 50856 148384 50862 148396
rect 185854 148384 185860 148396
rect 185912 148384 185918 148436
rect 407022 148384 407028 148436
rect 407080 148424 407086 148436
rect 525886 148424 525892 148436
rect 407080 148396 525892 148424
rect 407080 148384 407086 148396
rect 525886 148384 525892 148396
rect 525944 148384 525950 148436
rect 48314 148316 48320 148368
rect 48372 148356 48378 148368
rect 188798 148356 188804 148368
rect 48372 148328 188804 148356
rect 48372 148316 48378 148328
rect 188798 148316 188804 148328
rect 188856 148316 188862 148368
rect 410978 148316 410984 148368
rect 411036 148356 411042 148368
rect 531038 148356 531044 148368
rect 411036 148328 531044 148356
rect 411036 148316 411042 148328
rect 531038 148316 531044 148328
rect 531096 148316 531102 148368
rect 113450 148248 113456 148300
rect 113508 148288 113514 148300
rect 183094 148288 183100 148300
rect 113508 148260 183100 148288
rect 113508 148248 113514 148260
rect 183094 148248 183100 148260
rect 183152 148248 183158 148300
rect 406562 148248 406568 148300
rect 406620 148288 406626 148300
rect 465994 148288 466000 148300
rect 406620 148260 466000 148288
rect 406620 148248 406626 148260
rect 465994 148248 466000 148260
rect 466052 148248 466058 148300
rect 115842 148180 115848 148232
rect 115900 148220 115906 148232
rect 183002 148220 183008 148232
rect 115900 148192 183008 148220
rect 115900 148180 115906 148192
rect 183002 148180 183008 148192
rect 183060 148180 183066 148232
rect 406746 148180 406752 148232
rect 406804 148220 406810 148232
rect 463510 148220 463516 148232
rect 406804 148192 463516 148220
rect 406804 148180 406810 148192
rect 463510 148180 463516 148192
rect 463568 148180 463574 148232
rect 120902 148112 120908 148164
rect 120960 148152 120966 148164
rect 182818 148152 182824 148164
rect 120960 148124 182824 148152
rect 120960 148112 120966 148124
rect 182818 148112 182824 148124
rect 182876 148112 182882 148164
rect 17034 147840 17040 147892
rect 17092 147880 17098 147892
rect 19702 147880 19708 147892
rect 17092 147852 19708 147880
rect 17092 147840 17098 147852
rect 19702 147840 19708 147852
rect 19760 147840 19766 147892
rect 19978 147840 19984 147892
rect 20036 147880 20042 147892
rect 48222 147880 48228 147892
rect 20036 147852 48228 147880
rect 20036 147840 20042 147852
rect 48222 147840 48228 147852
rect 48280 147840 48286 147892
rect 48130 147812 48136 147824
rect 18708 147784 48136 147812
rect 18708 147756 18736 147784
rect 48130 147772 48136 147784
rect 48188 147772 48194 147824
rect 18138 147704 18144 147756
rect 18196 147744 18202 147756
rect 18690 147744 18696 147756
rect 18196 147716 18696 147744
rect 18196 147704 18202 147716
rect 18690 147704 18696 147716
rect 18748 147704 18754 147756
rect 58066 147744 58072 147756
rect 19260 147716 58072 147744
rect 19260 147688 19288 147716
rect 58066 147704 58072 147716
rect 58124 147744 58130 147756
rect 59354 147744 59360 147756
rect 58124 147716 59360 147744
rect 58124 147704 58130 147716
rect 59354 147704 59360 147716
rect 59412 147704 59418 147756
rect 18230 147636 18236 147688
rect 18288 147676 18294 147688
rect 19242 147676 19248 147688
rect 18288 147648 19248 147676
rect 18288 147636 18294 147648
rect 19242 147636 19248 147648
rect 19300 147636 19306 147688
rect 19702 147636 19708 147688
rect 19760 147676 19766 147688
rect 59538 147676 59544 147688
rect 19760 147648 59544 147676
rect 19760 147636 19766 147648
rect 59538 147636 59544 147648
rect 59596 147636 59602 147688
rect 19058 147568 19064 147620
rect 19116 147608 19122 147620
rect 36998 147608 37004 147620
rect 19116 147580 37004 147608
rect 19116 147568 19122 147580
rect 36998 147568 37004 147580
rect 37056 147568 37062 147620
rect 48222 147568 48228 147620
rect 48280 147608 48286 147620
rect 50154 147608 50160 147620
rect 48280 147580 50160 147608
rect 48280 147568 48286 147580
rect 50154 147568 50160 147580
rect 50212 147568 50218 147620
rect 63586 147568 63592 147620
rect 63644 147608 63650 147620
rect 189718 147608 189724 147620
rect 63644 147580 189724 147608
rect 63644 147568 63650 147580
rect 189718 147568 189724 147580
rect 189776 147568 189782 147620
rect 406470 147568 406476 147620
rect 406528 147608 406534 147620
rect 458358 147608 458364 147620
rect 406528 147580 458364 147608
rect 406528 147568 406534 147580
rect 458358 147568 458364 147580
rect 458416 147568 458422 147620
rect 459462 147568 459468 147620
rect 459520 147608 459526 147620
rect 478046 147608 478052 147620
rect 459520 147580 478052 147608
rect 459520 147568 459526 147580
rect 478046 147568 478052 147580
rect 478104 147568 478110 147620
rect 16114 147500 16120 147552
rect 16172 147540 16178 147552
rect 19334 147540 19340 147552
rect 16172 147512 19340 147540
rect 16172 147500 16178 147512
rect 19334 147500 19340 147512
rect 19392 147540 19398 147552
rect 20622 147540 20628 147552
rect 19392 147512 20628 147540
rect 19392 147500 19398 147512
rect 20622 147500 20628 147512
rect 20680 147500 20686 147552
rect 61654 147540 61660 147552
rect 45526 147512 61660 147540
rect 35894 147472 35900 147484
rect 18984 147444 35900 147472
rect 18984 147348 19012 147444
rect 35894 147432 35900 147444
rect 35952 147432 35958 147484
rect 19150 147364 19156 147416
rect 19208 147404 19214 147416
rect 38102 147404 38108 147416
rect 19208 147376 38108 147404
rect 19208 147364 19214 147376
rect 38102 147364 38108 147376
rect 38160 147364 38166 147416
rect 18598 147296 18604 147348
rect 18656 147336 18662 147348
rect 18966 147336 18972 147348
rect 18656 147308 18972 147336
rect 18656 147296 18662 147308
rect 18966 147296 18972 147308
rect 19024 147296 19030 147348
rect 19886 147296 19892 147348
rect 19944 147336 19950 147348
rect 43070 147336 43076 147348
rect 19944 147308 43076 147336
rect 19944 147296 19950 147308
rect 43070 147296 43076 147308
rect 43128 147336 43134 147348
rect 45526 147336 45554 147512
rect 61654 147500 61660 147512
rect 61712 147500 61718 147552
rect 66162 147500 66168 147552
rect 66220 147540 66226 147552
rect 180058 147540 180064 147552
rect 66220 147512 180064 147540
rect 66220 147500 66226 147512
rect 180058 147500 180064 147512
rect 180116 147500 180122 147552
rect 406654 147500 406660 147552
rect 406712 147540 406718 147552
rect 455966 147540 455972 147552
rect 406712 147512 455972 147540
rect 406712 147500 406718 147512
rect 455966 147500 455972 147512
rect 456024 147500 456030 147552
rect 458082 147500 458088 147552
rect 458140 147540 458146 147552
rect 476942 147540 476948 147552
rect 458140 147512 476948 147540
rect 458140 147500 458146 147512
rect 476942 147500 476948 147512
rect 477000 147500 477006 147552
rect 48130 147432 48136 147484
rect 48188 147472 48194 147484
rect 51442 147472 51448 147484
rect 48188 147444 51448 147472
rect 48188 147432 48194 147444
rect 51442 147432 51448 147444
rect 51500 147432 51506 147484
rect 59538 147432 59544 147484
rect 59596 147472 59602 147484
rect 78030 147472 78036 147484
rect 59596 147444 78036 147472
rect 59596 147432 59602 147444
rect 78030 147432 78036 147444
rect 78088 147432 78094 147484
rect 78490 147432 78496 147484
rect 78548 147472 78554 147484
rect 188430 147472 188436 147484
rect 78548 147444 188436 147472
rect 78548 147432 78554 147444
rect 188430 147432 188436 147444
rect 188488 147432 188494 147484
rect 409138 147432 409144 147484
rect 409196 147472 409202 147484
rect 453574 147472 453580 147484
rect 409196 147444 453580 147472
rect 409196 147432 409202 147444
rect 453574 147432 453580 147444
rect 453632 147432 453638 147484
rect 47670 147364 47676 147416
rect 47728 147404 47734 147416
rect 66346 147404 66352 147416
rect 47728 147376 66352 147404
rect 47728 147364 47734 147376
rect 66346 147364 66352 147376
rect 66404 147364 66410 147416
rect 70394 147364 70400 147416
rect 70452 147404 70458 147416
rect 75638 147404 75644 147416
rect 70452 147376 75644 147404
rect 70452 147364 70458 147376
rect 75638 147364 75644 147376
rect 75696 147364 75702 147416
rect 75822 147364 75828 147416
rect 75880 147404 75886 147416
rect 79134 147404 79140 147416
rect 75880 147376 79140 147404
rect 75880 147364 75886 147376
rect 79134 147364 79140 147376
rect 79192 147364 79198 147416
rect 81066 147364 81072 147416
rect 81124 147404 81130 147416
rect 188338 147404 188344 147416
rect 81124 147376 188344 147404
rect 81124 147364 81130 147376
rect 188338 147364 188344 147376
rect 188396 147364 188402 147416
rect 415118 147364 415124 147416
rect 415176 147404 415182 147416
rect 448238 147404 448244 147416
rect 415176 147376 448244 147404
rect 415176 147364 415182 147376
rect 448238 147364 448244 147376
rect 448296 147364 448302 147416
rect 43128 147308 45554 147336
rect 43128 147296 43134 147308
rect 59354 147296 59360 147348
rect 59412 147336 59418 147348
rect 76926 147336 76932 147348
rect 59412 147308 76932 147336
rect 59412 147296 59418 147308
rect 76926 147296 76932 147308
rect 76984 147296 76990 147348
rect 88242 147296 88248 147348
rect 88300 147336 88306 147348
rect 186038 147336 186044 147348
rect 88300 147308 186044 147336
rect 88300 147296 88306 147308
rect 186038 147296 186044 147308
rect 186096 147296 186102 147348
rect 418338 147296 418344 147348
rect 418396 147336 418402 147348
rect 450630 147336 450636 147348
rect 418396 147308 450636 147336
rect 418396 147296 418402 147308
rect 450630 147296 450636 147308
rect 450688 147296 450694 147348
rect 15654 147228 15660 147280
rect 15712 147268 15718 147280
rect 19242 147268 19248 147280
rect 15712 147240 19248 147268
rect 15712 147228 15718 147240
rect 19242 147228 19248 147240
rect 19300 147228 19306 147280
rect 19794 147228 19800 147280
rect 19852 147268 19858 147280
rect 44174 147268 44180 147280
rect 19852 147240 44180 147268
rect 19852 147228 19858 147240
rect 44174 147228 44180 147240
rect 44232 147268 44238 147280
rect 44726 147268 44732 147280
rect 44232 147240 44732 147268
rect 44232 147228 44238 147240
rect 44726 147228 44732 147240
rect 44784 147228 44790 147280
rect 46014 147228 46020 147280
rect 46072 147268 46078 147280
rect 46566 147268 46572 147280
rect 46072 147240 46572 147268
rect 46072 147228 46078 147240
rect 46566 147228 46572 147240
rect 46624 147268 46630 147280
rect 65150 147268 65156 147280
rect 46624 147240 65156 147268
rect 46624 147228 46630 147240
rect 65150 147228 65156 147240
rect 65208 147228 65214 147280
rect 91002 147228 91008 147280
rect 91060 147268 91066 147280
rect 185578 147268 185584 147280
rect 91060 147240 185584 147268
rect 91060 147228 91066 147240
rect 185578 147228 185584 147240
rect 185636 147228 185642 147280
rect 414658 147228 414664 147280
rect 414716 147268 414722 147280
rect 440234 147268 440240 147280
rect 414716 147240 440240 147268
rect 414716 147228 414722 147240
rect 440234 147228 440240 147240
rect 440292 147228 440298 147280
rect 15930 147160 15936 147212
rect 15988 147200 15994 147212
rect 16390 147200 16396 147212
rect 15988 147172 16396 147200
rect 15988 147160 15994 147172
rect 16390 147160 16396 147172
rect 16448 147200 16454 147212
rect 48682 147200 48688 147212
rect 16448 147172 48688 147200
rect 16448 147160 16454 147172
rect 48682 147160 48688 147172
rect 48740 147200 48746 147212
rect 67634 147200 67640 147212
rect 48740 147172 67640 147200
rect 48740 147160 48746 147172
rect 67634 147160 67640 147172
rect 67692 147160 67698 147212
rect 68278 147160 68284 147212
rect 68336 147200 68342 147212
rect 162210 147200 162216 147212
rect 68336 147172 162216 147200
rect 68336 147160 68342 147172
rect 162210 147160 162216 147172
rect 162268 147160 162274 147212
rect 418706 147160 418712 147212
rect 418764 147200 418770 147212
rect 419074 147200 419080 147212
rect 418764 147172 419080 147200
rect 418764 147160 418770 147172
rect 419074 147160 419080 147172
rect 419132 147200 419138 147212
rect 437014 147200 437020 147212
rect 419132 147172 437020 147200
rect 419132 147160 419138 147172
rect 437014 147160 437020 147172
rect 437072 147160 437078 147212
rect 18690 147092 18696 147144
rect 18748 147132 18754 147144
rect 19150 147132 19156 147144
rect 18748 147104 19156 147132
rect 18748 147092 18754 147104
rect 19150 147092 19156 147104
rect 19208 147092 19214 147144
rect 19702 147092 19708 147144
rect 19760 147132 19766 147144
rect 19886 147132 19892 147144
rect 19760 147104 19892 147132
rect 19760 147092 19766 147104
rect 19886 147092 19892 147104
rect 19944 147092 19950 147144
rect 21358 147092 21364 147144
rect 21416 147132 21422 147144
rect 54018 147132 54024 147144
rect 21416 147104 54024 147132
rect 21416 147092 21422 147104
rect 54018 147092 54024 147104
rect 54076 147092 54082 147144
rect 71222 147092 71228 147144
rect 71280 147132 71286 147144
rect 164050 147132 164056 147144
rect 71280 147104 164056 147132
rect 71280 147092 71286 147104
rect 164050 147092 164056 147104
rect 164108 147092 164114 147144
rect 419350 147092 419356 147144
rect 419408 147132 419414 147144
rect 439590 147132 439596 147144
rect 419408 147104 439596 147132
rect 419408 147092 419414 147104
rect 439590 147092 439596 147104
rect 439648 147092 439654 147144
rect 16022 147024 16028 147076
rect 16080 147064 16086 147076
rect 16482 147064 16488 147076
rect 16080 147036 16488 147064
rect 16080 147024 16086 147036
rect 16482 147024 16488 147036
rect 16540 147064 16546 147076
rect 52270 147064 52276 147076
rect 16540 147036 52276 147064
rect 16540 147024 16546 147036
rect 52270 147024 52276 147036
rect 52328 147064 52334 147076
rect 71038 147064 71044 147076
rect 52328 147036 71044 147064
rect 52328 147024 52334 147036
rect 71038 147024 71044 147036
rect 71096 147024 71102 147076
rect 95970 147024 95976 147076
rect 96028 147064 96034 147076
rect 185762 147064 185768 147076
rect 96028 147036 185768 147064
rect 96028 147024 96034 147036
rect 185762 147024 185768 147036
rect 185820 147024 185826 147076
rect 419626 147024 419632 147076
rect 419684 147064 419690 147076
rect 443086 147064 443092 147076
rect 419684 147036 443092 147064
rect 419684 147024 419690 147036
rect 443086 147024 443092 147036
rect 443144 147064 443150 147076
rect 461670 147064 461676 147076
rect 443144 147036 461676 147064
rect 443144 147024 443150 147036
rect 461670 147024 461676 147036
rect 461728 147024 461734 147076
rect 16298 146956 16304 147008
rect 16356 146996 16362 147008
rect 53374 146996 53380 147008
rect 16356 146968 53380 146996
rect 16356 146956 16362 146968
rect 53374 146956 53380 146968
rect 53432 146996 53438 147008
rect 72142 146996 72148 147008
rect 53432 146968 72148 146996
rect 53432 146956 53438 146968
rect 72142 146956 72148 146968
rect 72200 146956 72206 147008
rect 103514 146956 103520 147008
rect 103572 146996 103578 147008
rect 191098 146996 191104 147008
rect 103572 146968 191104 146996
rect 103572 146956 103578 146968
rect 191098 146956 191104 146968
rect 191156 146956 191162 147008
rect 418430 146956 418436 147008
rect 418488 146996 418494 147008
rect 419258 146996 419264 147008
rect 418488 146968 419264 146996
rect 418488 146956 418494 146968
rect 419258 146956 419264 146968
rect 419316 146996 419322 147008
rect 444190 146996 444196 147008
rect 419316 146968 444196 146996
rect 419316 146956 419322 146968
rect 444190 146956 444196 146968
rect 444248 146996 444254 147008
rect 462774 146996 462780 147008
rect 444248 146968 462780 146996
rect 444248 146956 444254 146968
rect 462774 146956 462780 146968
rect 462832 146956 462838 147008
rect 18874 146888 18880 146940
rect 18932 146928 18938 146940
rect 21358 146928 21364 146940
rect 18932 146900 21364 146928
rect 18932 146888 18938 146900
rect 21358 146888 21364 146900
rect 21416 146888 21422 146940
rect 56042 146928 56048 146940
rect 26206 146900 56048 146928
rect 18322 146820 18328 146872
rect 18380 146860 18386 146872
rect 26206 146860 26234 146900
rect 56042 146888 56048 146900
rect 56100 146928 56106 146940
rect 73706 146928 73712 146940
rect 56100 146900 73712 146928
rect 56100 146888 56106 146900
rect 73706 146888 73712 146900
rect 73764 146888 73770 146940
rect 100938 146888 100944 146940
rect 100996 146928 101002 146940
rect 182910 146928 182916 146940
rect 100996 146900 182916 146928
rect 100996 146888 101002 146900
rect 182910 146888 182916 146900
rect 182968 146888 182974 146940
rect 419718 146888 419724 146940
rect 419776 146928 419782 146940
rect 419902 146928 419908 146940
rect 419776 146900 419908 146928
rect 419776 146888 419782 146900
rect 419902 146888 419908 146900
rect 419960 146928 419966 146940
rect 454586 146928 454592 146940
rect 419960 146900 454592 146928
rect 419960 146888 419966 146900
rect 454586 146888 454592 146900
rect 454644 146928 454650 146940
rect 473354 146928 473360 146940
rect 454644 146900 473360 146928
rect 454644 146888 454650 146900
rect 473354 146888 473360 146900
rect 473412 146888 473418 146940
rect 18380 146832 26234 146860
rect 18380 146820 18386 146832
rect 50154 146820 50160 146872
rect 50212 146860 50218 146872
rect 68462 146860 68468 146872
rect 50212 146832 68468 146860
rect 50212 146820 50218 146832
rect 68462 146820 68468 146832
rect 68520 146820 68526 146872
rect 106090 146820 106096 146872
rect 106148 146860 106154 146872
rect 156598 146860 156604 146872
rect 106148 146832 156604 146860
rect 106148 146820 106154 146832
rect 156598 146820 156604 146832
rect 156656 146820 156662 146872
rect 418614 146820 418620 146872
rect 418672 146860 418678 146872
rect 419166 146860 419172 146872
rect 418672 146832 419172 146860
rect 418672 146820 418678 146832
rect 419166 146820 419172 146832
rect 419224 146860 419230 146872
rect 437934 146860 437940 146872
rect 419224 146832 437940 146860
rect 419224 146820 419230 146832
rect 437934 146820 437940 146832
rect 437992 146820 437998 146872
rect 445294 146820 445300 146872
rect 445352 146860 445358 146872
rect 463878 146860 463884 146872
rect 445352 146832 463884 146860
rect 445352 146820 445358 146832
rect 463878 146820 463884 146832
rect 463936 146820 463942 146872
rect 51442 146752 51448 146804
rect 51500 146792 51506 146804
rect 69750 146792 69756 146804
rect 51500 146764 69756 146792
rect 51500 146752 51506 146764
rect 69750 146752 69756 146764
rect 69808 146752 69814 146804
rect 108850 146752 108856 146804
rect 108908 146792 108914 146804
rect 158162 146792 158168 146804
rect 108908 146764 158168 146792
rect 108908 146752 108914 146764
rect 158162 146752 158168 146764
rect 158220 146752 158226 146804
rect 418890 146752 418896 146804
rect 418948 146792 418954 146804
rect 436094 146792 436100 146804
rect 418948 146764 436100 146792
rect 418948 146752 418954 146764
rect 436094 146752 436100 146764
rect 436152 146752 436158 146804
rect 447134 146752 447140 146804
rect 447192 146792 447198 146804
rect 466270 146792 466276 146804
rect 447192 146764 466276 146792
rect 447192 146752 447198 146764
rect 466270 146752 466276 146764
rect 466328 146752 466334 146804
rect 45278 146724 45284 146736
rect 42260 146696 45284 146724
rect 18782 146480 18788 146532
rect 18840 146520 18846 146532
rect 39574 146520 39580 146532
rect 18840 146492 39580 146520
rect 18840 146480 18846 146492
rect 39574 146480 39580 146492
rect 39632 146480 39638 146532
rect 18506 146412 18512 146464
rect 18564 146452 18570 146464
rect 19242 146452 19248 146464
rect 18564 146424 19248 146452
rect 18564 146412 18570 146424
rect 19242 146412 19248 146424
rect 19300 146452 19306 146464
rect 42260 146452 42288 146696
rect 45278 146684 45284 146696
rect 45336 146724 45342 146736
rect 63862 146724 63868 146736
rect 45336 146696 63868 146724
rect 45336 146684 45342 146696
rect 63862 146684 63868 146696
rect 63920 146684 63926 146736
rect 111610 146684 111616 146736
rect 111668 146724 111674 146736
rect 157978 146724 157984 146736
rect 111668 146696 157984 146724
rect 111668 146684 111674 146696
rect 157978 146684 157984 146696
rect 158036 146684 158042 146736
rect 430574 146684 430580 146736
rect 430632 146724 430638 146736
rect 438210 146724 438216 146736
rect 430632 146696 438216 146724
rect 430632 146684 430638 146696
rect 438210 146684 438216 146696
rect 438268 146684 438274 146736
rect 448514 146684 448520 146736
rect 448572 146724 448578 146736
rect 467558 146724 467564 146736
rect 448572 146696 467564 146724
rect 448572 146684 448578 146696
rect 467558 146684 467564 146696
rect 467616 146684 467622 146736
rect 44726 146616 44732 146668
rect 44784 146656 44790 146668
rect 62758 146656 62764 146668
rect 44784 146628 62764 146656
rect 44784 146616 44790 146628
rect 62758 146616 62764 146628
rect 62816 146616 62822 146668
rect 449894 146616 449900 146668
rect 449952 146656 449958 146668
rect 468662 146656 468668 146668
rect 449952 146628 468668 146656
rect 449952 146616 449958 146628
rect 468662 146616 468668 146628
rect 468720 146616 468726 146668
rect 54018 146548 54024 146600
rect 54076 146588 54082 146600
rect 73246 146588 73252 146600
rect 54076 146560 73252 146588
rect 54076 146548 54082 146560
rect 73246 146548 73252 146560
rect 73304 146548 73310 146600
rect 452470 146548 452476 146600
rect 452528 146588 452534 146600
rect 469766 146588 469772 146600
rect 452528 146560 469772 146588
rect 452528 146548 452534 146560
rect 469766 146548 469772 146560
rect 469824 146548 469830 146600
rect 452562 146480 452568 146532
rect 452620 146520 452626 146532
rect 471054 146520 471060 146532
rect 452620 146492 471060 146520
rect 452620 146480 452626 146492
rect 471054 146480 471060 146492
rect 471112 146480 471118 146532
rect 19300 146424 42288 146452
rect 19300 146412 19306 146424
rect 446398 146412 446404 146464
rect 446456 146452 446462 146464
rect 465166 146452 465172 146464
rect 446456 146424 465172 146452
rect 446456 146412 446462 146424
rect 465166 146412 465172 146424
rect 465224 146412 465230 146464
rect 15746 146344 15752 146396
rect 15804 146384 15810 146396
rect 18598 146384 18604 146396
rect 15804 146356 18604 146384
rect 15804 146344 15810 146356
rect 18598 146344 18604 146356
rect 18656 146384 18662 146396
rect 46014 146384 46020 146396
rect 18656 146356 46020 146384
rect 18656 146344 18662 146356
rect 46014 146344 46020 146356
rect 46072 146344 46078 146396
rect 472158 146384 472164 146396
rect 453960 146356 472164 146384
rect 20622 146276 20628 146328
rect 20680 146316 20686 146328
rect 47670 146316 47676 146328
rect 20680 146288 47676 146316
rect 20680 146276 20686 146288
rect 47670 146276 47676 146288
rect 47728 146276 47734 146328
rect 415762 146208 415768 146260
rect 415820 146248 415826 146260
rect 416314 146248 416320 146260
rect 415820 146220 416320 146248
rect 415820 146208 415826 146220
rect 416314 146208 416320 146220
rect 416372 146208 416378 146260
rect 417142 146208 417148 146260
rect 417200 146248 417206 146260
rect 417786 146248 417792 146260
rect 417200 146220 417792 146248
rect 417200 146208 417206 146220
rect 417786 146208 417792 146220
rect 417844 146208 417850 146260
rect 449894 146248 449900 146260
rect 418172 146220 449900 146248
rect 416332 146180 416360 146208
rect 418172 146180 418200 146220
rect 449894 146208 449900 146220
rect 449952 146208 449958 146260
rect 416332 146152 418200 146180
rect 419810 146140 419816 146192
rect 419868 146180 419874 146192
rect 453390 146180 453396 146192
rect 419868 146152 453396 146180
rect 419868 146140 419874 146152
rect 453390 146140 453396 146152
rect 453448 146180 453454 146192
rect 453960 146180 453988 146356
rect 472158 146344 472164 146356
rect 472216 146344 472222 146396
rect 456794 146276 456800 146328
rect 456852 146316 456858 146328
rect 474090 146316 474096 146328
rect 456852 146288 474096 146316
rect 456852 146276 456858 146288
rect 474090 146276 474096 146288
rect 474148 146276 474154 146328
rect 453448 146152 453988 146180
rect 453448 146140 453454 146152
rect 415670 146072 415676 146124
rect 415728 146112 415734 146124
rect 416682 146112 416688 146124
rect 415728 146084 416688 146112
rect 415728 146072 415734 146084
rect 416682 146072 416688 146084
rect 416740 146072 416746 146124
rect 419442 146072 419448 146124
rect 419500 146112 419506 146124
rect 452562 146112 452568 146124
rect 419500 146084 452568 146112
rect 419500 146072 419506 146084
rect 452562 146072 452568 146084
rect 452620 146072 452626 146124
rect 416700 146044 416728 146072
rect 448514 146044 448520 146056
rect 416700 146016 448520 146044
rect 448514 146004 448520 146016
rect 448572 146004 448578 146056
rect 419534 145936 419540 145988
rect 419592 145976 419598 145988
rect 419994 145976 420000 145988
rect 419592 145948 420000 145976
rect 419592 145936 419598 145948
rect 419994 145936 420000 145948
rect 420052 145976 420058 145988
rect 451274 145976 451280 145988
rect 420052 145948 451280 145976
rect 420052 145936 420058 145948
rect 451274 145936 451280 145948
rect 451332 145976 451338 145988
rect 452470 145976 452476 145988
rect 451332 145948 452476 145976
rect 451332 145936 451338 145948
rect 452470 145936 452476 145948
rect 452528 145936 452534 145988
rect 416498 145868 416504 145920
rect 416556 145908 416562 145920
rect 447134 145908 447140 145920
rect 416556 145880 447140 145908
rect 416556 145868 416562 145880
rect 447134 145868 447140 145880
rect 447192 145868 447198 145920
rect 417786 145800 417792 145852
rect 417844 145840 417850 145852
rect 445294 145840 445300 145852
rect 417844 145812 445300 145840
rect 417844 145800 417850 145812
rect 445294 145800 445300 145812
rect 445352 145800 445358 145852
rect 418982 145732 418988 145784
rect 419040 145772 419046 145784
rect 446398 145772 446404 145784
rect 419040 145744 446404 145772
rect 419040 145732 419046 145744
rect 446398 145732 446404 145744
rect 446456 145732 446462 145784
rect 531038 144848 531044 144900
rect 531096 144888 531102 144900
rect 536834 144888 536840 144900
rect 531096 144860 536840 144888
rect 531096 144848 531102 144860
rect 536834 144848 536840 144860
rect 536892 144848 536898 144900
rect 577590 139340 577596 139392
rect 577648 139380 577654 139392
rect 579614 139380 579620 139392
rect 577648 139352 579620 139380
rect 577648 139340 577654 139352
rect 579614 139340 579620 139352
rect 579672 139340 579678 139392
rect 536834 138660 536840 138712
rect 536892 138700 536898 138712
rect 556890 138700 556896 138712
rect 536892 138672 556896 138700
rect 536892 138660 536898 138672
rect 556890 138660 556896 138672
rect 556948 138660 556954 138712
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 167822 137952 167828 137964
rect 3568 137924 167828 137952
rect 3568 137912 3574 137924
rect 167822 137912 167828 137924
rect 167880 137912 167886 137964
rect 151262 136552 151268 136604
rect 151320 136592 151326 136604
rect 156690 136592 156696 136604
rect 151320 136564 156696 136592
rect 151320 136552 151326 136564
rect 156690 136552 156696 136564
rect 156748 136552 156754 136604
rect 551922 136552 551928 136604
rect 551980 136592 551986 136604
rect 556798 136592 556804 136604
rect 551980 136564 556804 136592
rect 551980 136552 551986 136564
rect 556798 136552 556804 136564
rect 556856 136552 556862 136604
rect 418522 135192 418528 135244
rect 418580 135232 418586 135244
rect 456794 135232 456800 135244
rect 418580 135204 456800 135232
rect 418580 135192 418586 135204
rect 456794 135192 456800 135204
rect 456852 135192 456858 135244
rect 187510 134648 187516 134700
rect 187568 134688 187574 134700
rect 580442 134688 580448 134700
rect 187568 134660 580448 134688
rect 187568 134648 187574 134660
rect 580442 134648 580448 134660
rect 580500 134648 580506 134700
rect 187602 134580 187608 134632
rect 187660 134620 187666 134632
rect 580902 134620 580908 134632
rect 187660 134592 580908 134620
rect 187660 134580 187666 134592
rect 580902 134580 580908 134592
rect 580960 134580 580966 134632
rect 187418 134512 187424 134564
rect 187476 134552 187482 134564
rect 580350 134552 580356 134564
rect 187476 134524 580356 134552
rect 187476 134512 187482 134524
rect 580350 134512 580356 134524
rect 580408 134512 580414 134564
rect 417326 134376 417332 134428
rect 417384 134416 417390 134428
rect 418522 134416 418528 134428
rect 417384 134388 418528 134416
rect 417384 134376 417390 134388
rect 418522 134376 418528 134388
rect 418580 134376 418586 134428
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 14734 111772 14740 111784
rect 3200 111744 14740 111772
rect 3200 111732 3206 111744
rect 14734 111732 14740 111744
rect 14792 111732 14798 111784
rect 556890 110372 556896 110424
rect 556948 110412 556954 110424
rect 559558 110412 559564 110424
rect 556948 110384 559564 110412
rect 556948 110372 556954 110384
rect 559558 110372 559564 110384
rect 559616 110372 559622 110424
rect 577498 100648 577504 100700
rect 577556 100688 577562 100700
rect 579706 100688 579712 100700
rect 577556 100660 579712 100688
rect 577556 100648 577562 100660
rect 579706 100648 579712 100660
rect 579764 100648 579770 100700
rect 559558 98948 559564 99000
rect 559616 98988 559622 99000
rect 565078 98988 565084 99000
rect 559616 98960 565084 98988
rect 559616 98948 559622 98960
rect 565078 98948 565084 98960
rect 565136 98948 565142 99000
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 14642 97968 14648 97980
rect 3568 97940 14648 97968
rect 3568 97928 3574 97940
rect 14642 97928 14648 97940
rect 14700 97928 14706 97980
rect 565078 91740 565084 91792
rect 565136 91780 565142 91792
rect 569954 91780 569960 91792
rect 565136 91752 569960 91780
rect 565136 91740 565142 91752
rect 569954 91740 569960 91752
rect 570012 91740 570018 91792
rect 161474 88952 161480 89004
rect 161532 88992 161538 89004
rect 211154 88992 211160 89004
rect 161532 88964 211160 88992
rect 161532 88952 161538 88964
rect 211154 88952 211160 88964
rect 211212 88952 211218 89004
rect 269114 88952 269120 89004
rect 269172 88992 269178 89004
rect 309778 88992 309784 89004
rect 269172 88964 309784 88992
rect 269172 88952 269178 88964
rect 309778 88952 309784 88964
rect 309836 88952 309842 89004
rect 267734 87592 267740 87644
rect 267792 87632 267798 87644
rect 305638 87632 305644 87644
rect 267792 87604 305644 87632
rect 267792 87592 267798 87604
rect 305638 87592 305644 87604
rect 305696 87592 305702 87644
rect 233878 87320 233884 87372
rect 233936 87360 233942 87372
rect 234614 87360 234620 87372
rect 233936 87332 234620 87360
rect 233936 87320 233942 87332
rect 234614 87320 234620 87332
rect 234672 87320 234678 87372
rect 190454 86232 190460 86284
rect 190512 86272 190518 86284
rect 222194 86272 222200 86284
rect 190512 86244 222200 86272
rect 190512 86232 190518 86244
rect 222194 86232 222200 86244
rect 222252 86232 222258 86284
rect 302878 86232 302884 86284
rect 302936 86272 302942 86284
rect 389174 86272 389180 86284
rect 302936 86244 389180 86272
rect 302936 86232 302942 86244
rect 389174 86232 389180 86244
rect 389232 86232 389238 86284
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 14550 85524 14556 85536
rect 3568 85496 14556 85524
rect 3568 85484 3574 85496
rect 14550 85484 14556 85496
rect 14608 85484 14614 85536
rect 569954 85484 569960 85536
rect 570012 85524 570018 85536
rect 573358 85524 573364 85536
rect 570012 85496 573364 85524
rect 570012 85484 570018 85496
rect 573358 85484 573364 85496
rect 573416 85484 573422 85536
rect 573358 73108 573364 73160
rect 573416 73148 573422 73160
rect 580166 73148 580172 73160
rect 573416 73120 580172 73148
rect 573416 73108 573422 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 14458 71720 14464 71732
rect 3568 71692 14464 71720
rect 3568 71680 3574 71692
rect 14458 71680 14464 71692
rect 14516 71680 14522 71732
rect 393958 59304 393964 59356
rect 394016 59344 394022 59356
rect 416774 59344 416780 59356
rect 394016 59316 416780 59344
rect 394016 59304 394022 59316
rect 416774 59304 416780 59316
rect 416832 59304 416838 59356
rect 418706 49920 418712 49972
rect 418764 49960 418770 49972
rect 456978 49960 456984 49972
rect 418764 49932 456984 49960
rect 418764 49920 418770 49932
rect 456978 49920 456984 49932
rect 457036 49920 457042 49972
rect 16298 49852 16304 49904
rect 16356 49892 16362 49904
rect 53466 49892 53472 49904
rect 16356 49864 53472 49892
rect 16356 49852 16362 49864
rect 53466 49852 53472 49864
rect 53524 49852 53530 49904
rect 417694 49852 417700 49904
rect 417752 49892 417758 49904
rect 458082 49892 458088 49904
rect 417752 49864 458088 49892
rect 417752 49852 417758 49864
rect 458082 49852 458088 49864
rect 458140 49852 458146 49904
rect 17034 49784 17040 49836
rect 17092 49824 17098 49836
rect 59538 49824 59544 49836
rect 17092 49796 59544 49824
rect 17092 49784 17098 49796
rect 59538 49784 59544 49796
rect 59596 49784 59602 49836
rect 408310 49784 408316 49836
rect 408368 49824 408374 49836
rect 478506 49824 478512 49836
rect 408368 49796 478512 49824
rect 408368 49784 408374 49796
rect 478506 49784 478512 49796
rect 478564 49784 478570 49836
rect 15102 49716 15108 49768
rect 15160 49756 15166 49768
rect 60642 49756 60648 49768
rect 15160 49728 60648 49756
rect 15160 49716 15166 49728
rect 60642 49716 60648 49728
rect 60700 49716 60706 49768
rect 408034 49716 408040 49768
rect 408092 49756 408098 49768
rect 480898 49756 480904 49768
rect 408092 49728 480904 49756
rect 408092 49716 408098 49728
rect 480898 49716 480904 49728
rect 480956 49716 480962 49768
rect 95878 49648 95884 49700
rect 95936 49688 95942 49700
rect 166626 49688 166632 49700
rect 95936 49660 166632 49688
rect 95936 49648 95942 49660
rect 166626 49648 166632 49660
rect 166684 49648 166690 49700
rect 407850 49648 407856 49700
rect 407908 49688 407914 49700
rect 495894 49688 495900 49700
rect 407908 49660 495900 49688
rect 407908 49648 407914 49660
rect 495894 49648 495900 49660
rect 495952 49648 495958 49700
rect 91002 49580 91008 49632
rect 91060 49620 91066 49632
rect 166442 49620 166448 49632
rect 91060 49592 166448 49620
rect 91060 49580 91066 49592
rect 166442 49580 166448 49592
rect 166500 49580 166506 49632
rect 413554 49580 413560 49632
rect 413612 49620 413618 49632
rect 503530 49620 503536 49632
rect 413612 49592 503536 49620
rect 413612 49580 413618 49592
rect 503530 49580 503536 49592
rect 503588 49580 503594 49632
rect 88242 49512 88248 49564
rect 88300 49552 88306 49564
rect 166534 49552 166540 49564
rect 88300 49524 166540 49552
rect 88300 49512 88306 49524
rect 166534 49512 166540 49524
rect 166592 49512 166598 49564
rect 410794 49512 410800 49564
rect 410852 49552 410858 49564
rect 500954 49552 500960 49564
rect 410852 49524 500960 49552
rect 410852 49512 410858 49524
rect 500954 49512 500960 49524
rect 501012 49512 501018 49564
rect 86034 49444 86040 49496
rect 86092 49484 86098 49496
rect 166810 49484 166816 49496
rect 86092 49456 166816 49484
rect 86092 49444 86098 49456
rect 166810 49444 166816 49456
rect 166868 49444 166874 49496
rect 406378 49444 406384 49496
rect 406436 49484 406442 49496
rect 498470 49484 498476 49496
rect 406436 49456 498476 49484
rect 406436 49444 406442 49456
rect 498470 49444 498476 49456
rect 498528 49444 498534 49496
rect 83550 49376 83556 49428
rect 83608 49416 83614 49428
rect 166350 49416 166356 49428
rect 83608 49388 166356 49416
rect 83608 49376 83614 49388
rect 166350 49376 166356 49388
rect 166408 49376 166414 49428
rect 410886 49376 410892 49428
rect 410944 49416 410950 49428
rect 505922 49416 505928 49428
rect 410944 49388 505928 49416
rect 410944 49376 410950 49388
rect 505922 49376 505928 49388
rect 505980 49376 505986 49428
rect 80974 49308 80980 49360
rect 81032 49348 81038 49360
rect 166718 49348 166724 49360
rect 81032 49320 166724 49348
rect 81032 49308 81038 49320
rect 166718 49308 166724 49320
rect 166776 49308 166782 49360
rect 413646 49308 413652 49360
rect 413704 49348 413710 49360
rect 508498 49348 508504 49360
rect 413704 49320 508504 49348
rect 413704 49308 413710 49320
rect 508498 49308 508504 49320
rect 508556 49308 508562 49360
rect 58526 49240 58532 49292
rect 58584 49280 58590 49292
rect 159634 49280 159640 49292
rect 58584 49252 159640 49280
rect 58584 49240 58590 49252
rect 159634 49240 159640 49252
rect 159692 49240 159698 49292
rect 413462 49240 413468 49292
rect 413520 49280 413526 49292
rect 510982 49280 510988 49292
rect 413520 49252 510988 49280
rect 413520 49240 413526 49252
rect 510982 49240 510988 49252
rect 511040 49240 511046 49292
rect 56042 49172 56048 49224
rect 56100 49212 56106 49224
rect 159726 49212 159732 49224
rect 56100 49184 159732 49212
rect 56100 49172 56106 49184
rect 159726 49172 159732 49184
rect 159784 49172 159790 49224
rect 416130 49172 416136 49224
rect 416188 49212 416194 49224
rect 515858 49212 515864 49224
rect 416188 49184 515864 49212
rect 416188 49172 416194 49184
rect 515858 49172 515864 49184
rect 515916 49172 515922 49224
rect 53650 49104 53656 49156
rect 53708 49144 53714 49156
rect 161198 49144 161204 49156
rect 53708 49116 161204 49144
rect 53708 49104 53714 49116
rect 161198 49104 161204 49116
rect 161256 49104 161262 49156
rect 413370 49104 413376 49156
rect 413428 49144 413434 49156
rect 513374 49144 513380 49156
rect 413428 49116 513380 49144
rect 413428 49104 413434 49116
rect 513374 49104 513380 49116
rect 513432 49104 513438 49156
rect 50798 49036 50804 49088
rect 50856 49076 50862 49088
rect 163866 49076 163872 49088
rect 50856 49048 163872 49076
rect 50856 49036 50862 49048
rect 163866 49036 163872 49048
rect 163924 49036 163930 49088
rect 411898 49036 411904 49088
rect 411956 49076 411962 49088
rect 520918 49076 520924 49088
rect 411956 49048 520924 49076
rect 411956 49036 411962 49048
rect 520918 49036 520924 49048
rect 520976 49036 520982 49088
rect 48314 48968 48320 49020
rect 48372 49008 48378 49020
rect 169294 49008 169300 49020
rect 48372 48980 169300 49008
rect 48372 48968 48378 48980
rect 169294 48968 169300 48980
rect 169352 48968 169358 49020
rect 416590 48968 416596 49020
rect 416648 49008 416654 49020
rect 525886 49008 525892 49020
rect 416648 48980 525892 49008
rect 416648 48968 416654 48980
rect 525886 48968 525892 48980
rect 525944 48968 525950 49020
rect 98546 48900 98552 48952
rect 98604 48940 98610 48952
rect 163682 48940 163688 48952
rect 98604 48912 163688 48940
rect 98604 48900 98610 48912
rect 163682 48900 163688 48912
rect 163740 48900 163746 48952
rect 410610 48900 410616 48952
rect 410668 48940 410674 48952
rect 493410 48940 493416 48952
rect 410668 48912 493416 48940
rect 410668 48900 410674 48912
rect 493410 48900 493416 48912
rect 493468 48900 493474 48952
rect 103514 48832 103520 48884
rect 103572 48872 103578 48884
rect 163958 48872 163964 48884
rect 103572 48844 163964 48872
rect 103572 48832 103578 48844
rect 163958 48832 163964 48844
rect 164016 48832 164022 48884
rect 407942 48832 407948 48884
rect 408000 48872 408006 48884
rect 488258 48872 488264 48884
rect 408000 48844 488264 48872
rect 408000 48832 408006 48844
rect 488258 48832 488264 48844
rect 488316 48832 488322 48884
rect 105998 48764 106004 48816
rect 106056 48804 106062 48816
rect 163774 48804 163780 48816
rect 106056 48776 163780 48804
rect 106056 48764 106062 48776
rect 163774 48764 163780 48776
rect 163832 48764 163838 48816
rect 418798 48764 418804 48816
rect 418856 48804 418862 48816
rect 459922 48804 459928 48816
rect 418856 48776 459928 48804
rect 418856 48764 418862 48776
rect 459922 48764 459928 48776
rect 459980 48764 459986 48816
rect 19058 48220 19064 48272
rect 19116 48260 19122 48272
rect 36814 48260 36820 48272
rect 19116 48232 36820 48260
rect 19116 48220 19122 48232
rect 36814 48220 36820 48232
rect 36872 48220 36878 48272
rect 59538 48220 59544 48272
rect 59596 48260 59602 48272
rect 78030 48260 78036 48272
rect 59596 48232 78036 48260
rect 59596 48220 59602 48232
rect 78030 48220 78036 48232
rect 78088 48220 78094 48272
rect 125962 48220 125968 48272
rect 126020 48260 126026 48272
rect 388070 48260 388076 48272
rect 126020 48232 388076 48260
rect 126020 48220 126026 48232
rect 388070 48220 388076 48232
rect 388128 48220 388134 48272
rect 416038 48220 416044 48272
rect 416096 48260 416102 48272
rect 458358 48260 458364 48272
rect 416096 48232 458364 48260
rect 416096 48220 416102 48232
rect 458358 48220 458364 48232
rect 458416 48220 458422 48272
rect 459462 48220 459468 48272
rect 459520 48260 459526 48272
rect 478046 48260 478052 48272
rect 459520 48232 478052 48260
rect 459520 48220 459526 48232
rect 478046 48220 478052 48232
rect 478104 48220 478110 48272
rect 19610 48152 19616 48204
rect 19668 48192 19674 48204
rect 57054 48192 57060 48204
rect 19668 48164 57060 48192
rect 19668 48152 19674 48164
rect 57054 48152 57060 48164
rect 57112 48152 57118 48204
rect 61194 48152 61200 48204
rect 61252 48192 61258 48204
rect 159358 48192 159364 48204
rect 61252 48164 159364 48192
rect 61252 48152 61258 48164
rect 159358 48152 159364 48164
rect 159416 48152 159422 48204
rect 405090 48152 405096 48204
rect 405148 48192 405154 48204
rect 448238 48192 448244 48204
rect 405148 48164 448244 48192
rect 405148 48152 405154 48164
rect 448238 48152 448244 48164
rect 448296 48152 448302 48204
rect 458082 48152 458088 48204
rect 458140 48192 458146 48204
rect 476942 48192 476948 48204
rect 458140 48164 476948 48192
rect 458140 48152 458146 48164
rect 476942 48152 476948 48164
rect 477000 48152 477006 48204
rect 18414 48084 18420 48136
rect 18472 48124 18478 48136
rect 55858 48124 55864 48136
rect 18472 48096 55864 48124
rect 18472 48084 18478 48096
rect 55858 48084 55864 48096
rect 55916 48124 55922 48136
rect 56502 48124 56508 48136
rect 55916 48096 56508 48124
rect 55916 48084 55922 48096
rect 56502 48084 56508 48096
rect 56560 48084 56566 48136
rect 65978 48084 65984 48136
rect 66036 48124 66042 48136
rect 161106 48124 161112 48136
rect 66036 48096 161112 48124
rect 66036 48084 66042 48096
rect 161106 48084 161112 48096
rect 161164 48084 161170 48136
rect 413278 48084 413284 48136
rect 413336 48124 413342 48136
rect 453574 48124 453580 48136
rect 413336 48096 453580 48124
rect 413336 48084 413342 48096
rect 453574 48084 453580 48096
rect 453632 48084 453638 48136
rect 469122 48084 469128 48136
rect 469180 48124 469186 48136
rect 475654 48124 475660 48136
rect 469180 48096 475660 48124
rect 469180 48084 469186 48096
rect 475654 48084 475660 48096
rect 475712 48084 475718 48136
rect 18874 48016 18880 48068
rect 18932 48056 18938 48068
rect 18932 48028 52040 48056
rect 18932 48016 18938 48028
rect 16482 47948 16488 48000
rect 16540 47988 16546 48000
rect 16540 47960 51672 47988
rect 16540 47948 16546 47960
rect 16390 47880 16396 47932
rect 16448 47920 16454 47932
rect 48682 47920 48688 47932
rect 16448 47892 48688 47920
rect 16448 47880 16454 47892
rect 48682 47880 48688 47892
rect 48740 47920 48746 47932
rect 48740 47892 51580 47920
rect 48740 47880 48746 47892
rect 18138 47812 18144 47864
rect 18196 47852 18202 47864
rect 51442 47852 51448 47864
rect 18196 47824 51448 47852
rect 18196 47812 18202 47824
rect 51442 47812 51448 47824
rect 51500 47812 51506 47864
rect 19978 47744 19984 47796
rect 20036 47784 20042 47796
rect 49694 47784 49700 47796
rect 20036 47756 49700 47784
rect 20036 47744 20042 47756
rect 49694 47744 49700 47756
rect 49752 47744 49758 47796
rect 19334 47676 19340 47728
rect 19392 47716 19398 47728
rect 47578 47716 47584 47728
rect 19392 47688 47584 47716
rect 19392 47676 19398 47688
rect 47578 47676 47584 47688
rect 47636 47716 47642 47728
rect 48222 47716 48228 47728
rect 47636 47688 48228 47716
rect 47636 47676 47642 47688
rect 48222 47676 48228 47688
rect 48280 47676 48286 47728
rect 51552 47716 51580 47892
rect 51644 47784 51672 47960
rect 52012 47920 52040 48028
rect 63954 48016 63960 48068
rect 64012 48056 64018 48068
rect 159542 48056 159548 48068
rect 64012 48028 159548 48056
rect 64012 48016 64018 48028
rect 159542 48016 159548 48028
rect 159600 48016 159606 48068
rect 410518 48016 410524 48068
rect 410576 48056 410582 48068
rect 450630 48056 450636 48068
rect 410576 48028 450636 48056
rect 410576 48016 410582 48028
rect 450630 48016 450636 48028
rect 450688 48016 450694 48068
rect 53466 47948 53472 48000
rect 53524 47988 53530 48000
rect 71774 47988 71780 48000
rect 53524 47960 71780 47988
rect 53524 47948 53530 47960
rect 71774 47948 71780 47960
rect 71832 47948 71838 48000
rect 73798 47948 73804 48000
rect 73856 47988 73862 48000
rect 169110 47988 169116 48000
rect 73856 47960 169116 47988
rect 73856 47948 73862 47960
rect 169110 47948 169116 47960
rect 169168 47948 169174 48000
rect 417326 47948 417332 48000
rect 417384 47988 417390 48000
rect 455874 47988 455880 48000
rect 417384 47960 455880 47988
rect 417384 47948 417390 47960
rect 455874 47948 455880 47960
rect 455932 47988 455938 48000
rect 474366 47988 474372 48000
rect 455932 47960 474372 47988
rect 455932 47948 455938 47960
rect 474366 47948 474372 47960
rect 474424 47948 474430 48000
rect 54570 47920 54576 47932
rect 52012 47892 54576 47920
rect 54570 47880 54576 47892
rect 54628 47920 54634 47932
rect 73246 47920 73252 47932
rect 54628 47892 73252 47920
rect 54628 47880 54634 47892
rect 73246 47880 73252 47892
rect 73304 47880 73310 47932
rect 76098 47880 76104 47932
rect 76156 47920 76162 47932
rect 169202 47920 169208 47932
rect 76156 47892 169208 47920
rect 76156 47880 76162 47892
rect 169202 47880 169208 47892
rect 169260 47880 169266 47932
rect 419718 47880 419724 47932
rect 419776 47920 419782 47932
rect 454586 47920 454592 47932
rect 419776 47892 454592 47920
rect 419776 47880 419782 47892
rect 454586 47880 454592 47892
rect 454644 47920 454650 47932
rect 454644 47892 465764 47920
rect 454644 47880 454650 47892
rect 68370 47812 68376 47864
rect 68428 47852 68434 47864
rect 159450 47852 159456 47864
rect 68428 47824 159456 47852
rect 68428 47812 68434 47824
rect 159450 47812 159456 47824
rect 159508 47812 159514 47864
rect 419258 47812 419264 47864
rect 419316 47852 419322 47864
rect 444282 47852 444288 47864
rect 419316 47824 444288 47852
rect 419316 47812 419322 47824
rect 444282 47812 444288 47824
rect 444340 47812 444346 47864
rect 52362 47784 52368 47796
rect 51644 47756 52368 47784
rect 52362 47744 52368 47756
rect 52420 47784 52426 47796
rect 71038 47784 71044 47796
rect 52420 47756 71044 47784
rect 52420 47744 52426 47756
rect 71038 47744 71044 47756
rect 71096 47744 71102 47796
rect 71130 47744 71136 47796
rect 71188 47784 71194 47796
rect 162118 47784 162124 47796
rect 71188 47756 162124 47784
rect 71188 47744 71194 47756
rect 162118 47744 162124 47756
rect 162176 47744 162182 47796
rect 419626 47744 419632 47796
rect 419684 47784 419690 47796
rect 419684 47756 441614 47784
rect 419684 47744 419690 47756
rect 67634 47716 67640 47728
rect 51552 47688 67640 47716
rect 67634 47676 67640 47688
rect 67692 47676 67698 47728
rect 78490 47676 78496 47728
rect 78548 47716 78554 47728
rect 169018 47716 169024 47728
rect 78548 47688 169024 47716
rect 78548 47676 78554 47688
rect 169018 47676 169024 47688
rect 169076 47676 169082 47728
rect 419350 47676 419356 47728
rect 419408 47716 419414 47728
rect 439590 47716 439596 47728
rect 419408 47688 439596 47716
rect 419408 47676 419414 47688
rect 439590 47676 439596 47688
rect 439648 47676 439654 47728
rect 441586 47716 441614 47756
rect 443086 47716 443092 47728
rect 441586 47688 443092 47716
rect 443086 47676 443092 47688
rect 443144 47716 443150 47728
rect 461670 47716 461676 47728
rect 443144 47688 461676 47716
rect 443144 47676 443150 47688
rect 461670 47676 461676 47688
rect 461728 47676 461734 47728
rect 18598 47608 18604 47660
rect 18656 47648 18662 47660
rect 46566 47648 46572 47660
rect 18656 47620 46572 47648
rect 18656 47608 18662 47620
rect 46566 47608 46572 47620
rect 46624 47648 46630 47660
rect 65058 47648 65064 47660
rect 46624 47620 65064 47648
rect 46624 47608 46630 47620
rect 65058 47608 65064 47620
rect 65116 47608 65122 47660
rect 93578 47608 93584 47660
rect 93636 47648 93642 47660
rect 166258 47648 166264 47660
rect 93636 47620 166264 47648
rect 93636 47608 93642 47620
rect 166258 47608 166264 47620
rect 166316 47608 166322 47660
rect 419166 47608 419172 47660
rect 419224 47648 419230 47660
rect 438118 47648 438124 47660
rect 419224 47620 438124 47648
rect 419224 47608 419230 47620
rect 438118 47608 438124 47620
rect 438176 47608 438182 47660
rect 444282 47608 444288 47660
rect 444340 47648 444346 47660
rect 462774 47648 462780 47660
rect 444340 47620 462780 47648
rect 444340 47608 444346 47620
rect 462774 47608 462780 47620
rect 462832 47608 462838 47660
rect 18506 47540 18512 47592
rect 18564 47580 18570 47592
rect 45370 47580 45376 47592
rect 18564 47552 45376 47580
rect 18564 47540 18570 47552
rect 45370 47540 45376 47552
rect 45428 47580 45434 47592
rect 45428 47552 45554 47580
rect 45428 47540 45434 47552
rect 19794 47472 19800 47524
rect 19852 47512 19858 47524
rect 44174 47512 44180 47524
rect 19852 47484 44180 47512
rect 19852 47472 19858 47484
rect 44174 47472 44180 47484
rect 44232 47472 44238 47524
rect 45526 47512 45554 47552
rect 48222 47540 48228 47592
rect 48280 47580 48286 47592
rect 66254 47580 66260 47592
rect 48280 47552 66260 47580
rect 48280 47540 48286 47552
rect 66254 47540 66260 47552
rect 66312 47540 66318 47592
rect 100938 47540 100944 47592
rect 100996 47580 101002 47592
rect 163590 47580 163596 47592
rect 100996 47552 163596 47580
rect 100996 47540 101002 47552
rect 163590 47540 163596 47552
rect 163648 47540 163654 47592
rect 418890 47540 418896 47592
rect 418948 47580 418954 47592
rect 436094 47580 436100 47592
rect 418948 47552 436100 47580
rect 418948 47540 418954 47552
rect 436094 47540 436100 47552
rect 436152 47540 436158 47592
rect 465736 47580 465764 47892
rect 473354 47580 473360 47592
rect 465736 47552 473360 47580
rect 473354 47540 473360 47552
rect 473412 47540 473418 47592
rect 63862 47512 63868 47524
rect 45526 47484 63868 47512
rect 63862 47472 63868 47484
rect 63920 47472 63926 47524
rect 111150 47472 111156 47524
rect 111208 47512 111214 47524
rect 160738 47512 160744 47524
rect 111208 47484 160744 47512
rect 111208 47472 111214 47484
rect 160738 47472 160744 47484
rect 160796 47472 160802 47524
rect 419074 47472 419080 47524
rect 419132 47512 419138 47524
rect 437014 47512 437020 47524
rect 419132 47484 437020 47512
rect 419132 47472 419138 47484
rect 437014 47472 437020 47484
rect 437072 47472 437078 47524
rect 19702 47404 19708 47456
rect 19760 47444 19766 47456
rect 43162 47444 43168 47456
rect 19760 47416 43168 47444
rect 19760 47404 19766 47416
rect 43162 47404 43168 47416
rect 43220 47444 43226 47456
rect 61378 47444 61384 47456
rect 43220 47416 61384 47444
rect 43220 47404 43226 47416
rect 61378 47404 61384 47416
rect 61436 47404 61442 47456
rect 115842 47404 115848 47456
rect 115900 47444 115906 47456
rect 160922 47444 160928 47456
rect 115900 47416 160928 47444
rect 115900 47404 115906 47416
rect 160922 47404 160928 47416
rect 160980 47404 160986 47456
rect 451274 47404 451280 47456
rect 451332 47444 451338 47456
rect 469214 47444 469220 47456
rect 451332 47416 469220 47444
rect 451332 47404 451338 47416
rect 469214 47404 469220 47416
rect 469272 47404 469278 47456
rect 44174 47336 44180 47388
rect 44232 47376 44238 47388
rect 62206 47376 62212 47388
rect 44232 47348 62212 47376
rect 44232 47336 44238 47348
rect 62206 47336 62212 47348
rect 62264 47336 62270 47388
rect 118602 47336 118608 47388
rect 118660 47376 118666 47388
rect 160830 47376 160836 47388
rect 118660 47348 160836 47376
rect 118660 47336 118666 47348
rect 160830 47336 160836 47348
rect 160888 47336 160894 47388
rect 449526 47336 449532 47388
rect 449584 47376 449590 47388
rect 467558 47376 467564 47388
rect 449584 47348 467564 47376
rect 449584 47336 449590 47348
rect 467558 47336 467564 47348
rect 467616 47336 467622 47388
rect 18230 47268 18236 47320
rect 18288 47308 18294 47320
rect 57974 47308 57980 47320
rect 18288 47280 57980 47308
rect 18288 47268 18294 47280
rect 57974 47268 57980 47280
rect 58032 47308 58038 47320
rect 76374 47308 76380 47320
rect 58032 47280 76380 47308
rect 58032 47268 58038 47280
rect 76374 47268 76380 47280
rect 76432 47268 76438 47320
rect 450446 47268 450452 47320
rect 450504 47308 450510 47320
rect 468662 47308 468668 47320
rect 450504 47280 468668 47308
rect 450504 47268 450510 47280
rect 468662 47268 468668 47280
rect 468720 47268 468726 47320
rect 50246 47200 50252 47252
rect 50304 47240 50310 47252
rect 68554 47240 68560 47252
rect 50304 47212 68560 47240
rect 50304 47200 50310 47212
rect 68554 47200 68560 47212
rect 68612 47200 68618 47252
rect 447502 47200 447508 47252
rect 447560 47240 447566 47252
rect 466270 47240 466276 47252
rect 447560 47212 466276 47240
rect 447560 47200 447566 47212
rect 466270 47200 466276 47212
rect 466328 47200 466334 47252
rect 56502 47132 56508 47184
rect 56560 47172 56566 47184
rect 74350 47172 74356 47184
rect 56560 47144 74356 47172
rect 56560 47132 56566 47144
rect 74350 47132 74356 47144
rect 74408 47132 74414 47184
rect 451274 47132 451280 47184
rect 451332 47172 451338 47184
rect 452286 47172 452292 47184
rect 451332 47144 452292 47172
rect 451332 47132 451338 47144
rect 452286 47132 452292 47144
rect 452344 47172 452350 47184
rect 471238 47172 471244 47184
rect 452344 47144 471244 47172
rect 452344 47132 452350 47144
rect 471238 47132 471244 47144
rect 471296 47132 471302 47184
rect 51442 47064 51448 47116
rect 51500 47104 51506 47116
rect 69750 47104 69756 47116
rect 51500 47076 69756 47104
rect 51500 47064 51506 47076
rect 69750 47064 69756 47076
rect 69808 47064 69814 47116
rect 445294 47064 445300 47116
rect 445352 47104 445358 47116
rect 463878 47104 463884 47116
rect 445352 47076 463884 47104
rect 445352 47064 445358 47076
rect 463878 47064 463884 47076
rect 463936 47064 463942 47116
rect 446398 46996 446404 47048
rect 446456 47036 446462 47048
rect 465166 47036 465172 47048
rect 446456 47008 465172 47036
rect 446456 46996 446462 47008
rect 465166 46996 465172 47008
rect 465224 46996 465230 47048
rect 453942 46928 453948 46980
rect 454000 46968 454006 46980
rect 472158 46968 472164 46980
rect 454000 46940 472164 46968
rect 454000 46928 454006 46940
rect 472158 46928 472164 46940
rect 472216 46928 472222 46980
rect 108850 46860 108856 46912
rect 108908 46900 108914 46912
rect 163498 46900 163504 46912
rect 108908 46872 163504 46900
rect 108908 46860 108914 46872
rect 163498 46860 163504 46872
rect 163556 46860 163562 46912
rect 190270 46860 190276 46912
rect 190328 46900 190334 46912
rect 580166 46900 580172 46912
rect 190328 46872 580172 46900
rect 190328 46860 190334 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 395338 46792 395344 46844
rect 395396 46832 395402 46844
rect 470870 46832 470876 46844
rect 395396 46804 470876 46832
rect 395396 46792 395402 46804
rect 470870 46792 470876 46804
rect 470928 46792 470934 46844
rect 395522 46724 395528 46776
rect 395580 46764 395586 46776
rect 468294 46764 468300 46776
rect 395580 46736 468300 46764
rect 395580 46724 395586 46736
rect 468294 46724 468300 46736
rect 468352 46724 468358 46776
rect 395430 46656 395436 46708
rect 395488 46696 395494 46708
rect 465902 46696 465908 46708
rect 395488 46668 465908 46696
rect 395488 46656 395494 46668
rect 465902 46656 465908 46668
rect 465960 46656 465966 46708
rect 403618 46588 403624 46640
rect 403676 46628 403682 46640
rect 463510 46628 463516 46640
rect 403676 46600 463516 46628
rect 403676 46588 403682 46600
rect 463510 46588 463516 46600
rect 463568 46588 463574 46640
rect 419810 46520 419816 46572
rect 419868 46560 419874 46572
rect 453942 46560 453948 46572
rect 419868 46532 453948 46560
rect 419868 46520 419874 46532
rect 453942 46520 453948 46532
rect 454000 46520 454006 46572
rect 418982 46452 418988 46504
rect 419040 46492 419046 46504
rect 446398 46492 446404 46504
rect 419040 46464 446404 46492
rect 419040 46452 419046 46464
rect 446398 46452 446404 46464
rect 446456 46452 446462 46504
rect 417786 46384 417792 46436
rect 417844 46424 417850 46436
rect 445294 46424 445300 46436
rect 417844 46396 445300 46424
rect 417844 46384 417850 46396
rect 445294 46384 445300 46396
rect 445352 46384 445358 46436
rect 133874 46180 133880 46232
rect 133932 46220 133938 46232
rect 199378 46220 199384 46232
rect 133932 46192 199384 46220
rect 133932 46180 133938 46192
rect 199378 46180 199384 46192
rect 199436 46180 199442 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 167730 45540 167736 45552
rect 3476 45512 167736 45540
rect 3476 45500 3482 45512
rect 167730 45500 167736 45512
rect 167788 45500 167794 45552
rect 416314 45500 416320 45552
rect 416372 45540 416378 45552
rect 450078 45540 450084 45552
rect 416372 45512 450084 45540
rect 416372 45500 416378 45512
rect 450078 45500 450084 45512
rect 450136 45500 450142 45552
rect 416682 45432 416688 45484
rect 416740 45472 416746 45484
rect 449526 45472 449532 45484
rect 416740 45444 449532 45472
rect 416740 45432 416746 45444
rect 449526 45432 449532 45444
rect 449584 45432 449590 45484
rect 419442 45364 419448 45416
rect 419500 45404 419506 45416
rect 451274 45404 451280 45416
rect 419500 45376 451280 45404
rect 419500 45364 419506 45376
rect 451274 45364 451280 45376
rect 451332 45364 451338 45416
rect 419994 45296 420000 45348
rect 420052 45336 420058 45348
rect 451366 45336 451372 45348
rect 420052 45308 451372 45336
rect 420052 45296 420058 45308
rect 451366 45296 451372 45308
rect 451424 45296 451430 45348
rect 416498 45228 416504 45280
rect 416556 45268 416562 45280
rect 447502 45268 447508 45280
rect 416556 45240 447508 45268
rect 416556 45228 416562 45240
rect 447502 45228 447508 45240
rect 447560 45228 447566 45280
rect 340874 44820 340880 44872
rect 340932 44860 340938 44872
rect 494698 44860 494704 44872
rect 340932 44832 494704 44860
rect 340932 44820 340938 44832
rect 494698 44820 494704 44832
rect 494756 44820 494762 44872
rect 336734 43392 336740 43444
rect 336792 43432 336798 43444
rect 483658 43432 483664 43444
rect 336792 43404 483664 43432
rect 336792 43392 336798 43404
rect 483658 43392 483664 43404
rect 483716 43392 483722 43444
rect 126974 42032 126980 42084
rect 127032 42072 127038 42084
rect 197446 42072 197452 42084
rect 127032 42044 197452 42072
rect 127032 42032 127038 42044
rect 197446 42032 197452 42044
rect 197504 42032 197510 42084
rect 347774 42032 347780 42084
rect 347832 42072 347838 42084
rect 512638 42072 512644 42084
rect 347832 42044 512644 42072
rect 347832 42032 347838 42044
rect 512638 42032 512644 42044
rect 512696 42032 512702 42084
rect 351914 40672 351920 40724
rect 351972 40712 351978 40724
rect 523034 40712 523040 40724
rect 351972 40684 523040 40712
rect 351972 40672 351978 40684
rect 523034 40672 523040 40684
rect 523092 40672 523098 40724
rect 125594 39312 125600 39364
rect 125652 39352 125658 39364
rect 194594 39352 194600 39364
rect 125652 39324 194600 39352
rect 125652 39312 125658 39324
rect 194594 39312 194600 39324
rect 194652 39312 194658 39364
rect 343634 39312 343640 39364
rect 343692 39352 343698 39364
rect 502334 39352 502340 39364
rect 343692 39324 502340 39352
rect 343692 39312 343698 39324
rect 502334 39312 502340 39324
rect 502392 39312 502398 39364
rect 316034 37884 316040 37936
rect 316092 37924 316098 37936
rect 431954 37924 431960 37936
rect 316092 37896 431960 37924
rect 316092 37884 316098 37896
rect 431954 37884 431960 37896
rect 432012 37884 432018 37936
rect 361574 36524 361580 36576
rect 361632 36564 361638 36576
rect 547874 36564 547880 36576
rect 361632 36536 547880 36564
rect 361632 36524 361638 36536
rect 547874 36524 547880 36536
rect 547932 36524 547938 36576
rect 313918 35164 313924 35216
rect 313976 35204 313982 35216
rect 420914 35204 420920 35216
rect 313976 35176 420920 35204
rect 313976 35164 313982 35176
rect 420914 35164 420920 35176
rect 420972 35164 420978 35216
rect 364334 33736 364340 33788
rect 364392 33776 364398 33788
rect 555418 33776 555424 33788
rect 364392 33748 555424 33776
rect 364392 33736 364398 33748
rect 555418 33736 555424 33748
rect 555476 33736 555482 33788
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 167638 33096 167644 33108
rect 3200 33068 167644 33096
rect 3200 33056 3206 33068
rect 167638 33056 167644 33068
rect 167696 33056 167702 33108
rect 335998 32376 336004 32428
rect 336056 32416 336062 32428
rect 473354 32416 473360 32428
rect 336056 32388 473360 32416
rect 336056 32376 336062 32388
rect 473354 32376 473360 32388
rect 473412 32376 473418 32428
rect 321554 31016 321560 31068
rect 321612 31056 321618 31068
rect 445754 31056 445760 31068
rect 321612 31028 445760 31056
rect 321612 31016 321618 31028
rect 445754 31016 445760 31028
rect 445812 31016 445818 31068
rect 320174 29588 320180 29640
rect 320232 29628 320238 29640
rect 441614 29628 441620 29640
rect 320232 29600 441620 29628
rect 320232 29588 320238 29600
rect 441614 29588 441620 29600
rect 441672 29588 441678 29640
rect 317414 28228 317420 28280
rect 317472 28268 317478 28280
rect 434714 28268 434720 28280
rect 317472 28240 434720 28268
rect 317472 28228 317478 28240
rect 434714 28228 434720 28240
rect 434772 28228 434778 28280
rect 329098 26868 329104 26920
rect 329156 26908 329162 26920
rect 456794 26908 456800 26920
rect 329156 26880 456800 26908
rect 329156 26868 329162 26880
rect 456794 26868 456800 26880
rect 456852 26868 456858 26920
rect 318794 25508 318800 25560
rect 318852 25548 318858 25560
rect 438854 25548 438860 25560
rect 318852 25520 438860 25548
rect 318852 25508 318858 25520
rect 438854 25508 438860 25520
rect 438912 25508 438918 25560
rect 211154 24080 211160 24132
rect 211212 24120 211218 24132
rect 230474 24120 230480 24132
rect 211212 24092 230480 24120
rect 211212 24080 211218 24092
rect 230474 24080 230480 24092
rect 230532 24080 230538 24132
rect 322934 24080 322940 24132
rect 322992 24120 322998 24132
rect 448514 24120 448520 24132
rect 322992 24092 448520 24120
rect 322992 24080 322998 24092
rect 448514 24080 448520 24092
rect 448572 24080 448578 24132
rect 314654 22720 314660 22772
rect 314712 22760 314718 22772
rect 427814 22760 427820 22772
rect 314712 22732 427820 22760
rect 314712 22720 314718 22732
rect 427814 22720 427820 22732
rect 427872 22720 427878 22772
rect 313274 21360 313280 21412
rect 313332 21400 313338 21412
rect 423674 21400 423680 21412
rect 313332 21372 423680 21400
rect 313332 21360 313338 21372
rect 423674 21360 423680 21372
rect 423732 21360 423738 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 170490 20652 170496 20664
rect 3476 20624 170496 20652
rect 3476 20612 3482 20624
rect 170490 20612 170496 20624
rect 170548 20612 170554 20664
rect 310514 17212 310520 17264
rect 310572 17252 310578 17264
rect 416774 17252 416780 17264
rect 310572 17224 416780 17252
rect 310572 17212 310578 17224
rect 416774 17212 416780 17224
rect 416832 17212 416838 17264
rect 298738 15852 298744 15904
rect 298796 15892 298802 15904
rect 364610 15892 364616 15904
rect 298796 15864 364616 15892
rect 298796 15852 298802 15864
rect 364610 15852 364616 15864
rect 364668 15852 364674 15904
rect 367094 15852 367100 15904
rect 367152 15892 367158 15904
rect 563054 15892 563060 15904
rect 367152 15864 563060 15892
rect 367152 15852 367158 15864
rect 563054 15852 563060 15864
rect 563112 15852 563118 15904
rect 273254 14424 273260 14476
rect 273312 14464 273318 14476
rect 322106 14464 322112 14476
rect 273312 14436 322112 14464
rect 273312 14424 273318 14436
rect 322106 14424 322112 14436
rect 322164 14424 322170 14476
rect 345014 14424 345020 14476
rect 345072 14464 345078 14476
rect 506474 14464 506480 14476
rect 345072 14436 506480 14464
rect 345072 14424 345078 14436
rect 506474 14424 506480 14436
rect 506532 14424 506538 14476
rect 346394 13064 346400 13116
rect 346452 13104 346458 13116
rect 508498 13104 508504 13116
rect 346452 13076 508504 13104
rect 346452 13064 346458 13076
rect 508498 13064 508504 13076
rect 508556 13064 508562 13116
rect 270494 11704 270500 11756
rect 270552 11744 270558 11756
rect 314654 11744 314660 11756
rect 270552 11716 314660 11744
rect 270552 11704 270558 11716
rect 314654 11704 314660 11716
rect 314712 11704 314718 11756
rect 342254 11704 342260 11756
rect 342312 11744 342318 11756
rect 498930 11744 498936 11756
rect 342312 11716 498936 11744
rect 342312 11704 342318 11716
rect 498930 11704 498936 11716
rect 498988 11704 498994 11756
rect 266354 10276 266360 10328
rect 266412 10316 266418 10328
rect 303890 10316 303896 10328
rect 266412 10288 303896 10316
rect 266412 10276 266418 10288
rect 303890 10276 303896 10288
rect 303948 10276 303954 10328
rect 339494 10276 339500 10328
rect 339552 10316 339558 10328
rect 492306 10316 492312 10328
rect 339552 10288 492312 10316
rect 339552 10276 339558 10288
rect 492306 10276 492312 10288
rect 492364 10276 492370 10328
rect 169570 8916 169576 8968
rect 169628 8956 169634 8968
rect 213914 8956 213920 8968
rect 169628 8928 213920 8956
rect 169628 8916 169634 8928
rect 213914 8916 213920 8928
rect 213972 8916 213978 8968
rect 262214 8916 262220 8968
rect 262272 8956 262278 8968
rect 291930 8956 291936 8968
rect 262272 8928 291936 8956
rect 262272 8916 262278 8928
rect 291930 8916 291936 8928
rect 291988 8916 291994 8968
rect 338114 8916 338120 8968
rect 338172 8956 338178 8968
rect 488810 8956 488816 8968
rect 338172 8928 488816 8956
rect 338172 8916 338178 8928
rect 488810 8916 488816 8928
rect 488868 8916 488874 8968
rect 263594 7624 263600 7676
rect 263652 7664 263658 7676
rect 294046 7664 294052 7676
rect 263652 7636 294052 7664
rect 263652 7624 263658 7636
rect 294046 7624 294052 7636
rect 294104 7624 294110 7676
rect 130562 7556 130568 7608
rect 130620 7596 130626 7608
rect 198734 7596 198740 7608
rect 130620 7568 198740 7596
rect 130620 7556 130626 7568
rect 198734 7556 198740 7568
rect 198792 7556 198798 7608
rect 201494 7556 201500 7608
rect 201552 7596 201558 7608
rect 226334 7596 226340 7608
rect 201552 7568 226340 7596
rect 201552 7556 201558 7568
rect 226334 7556 226340 7568
rect 226392 7556 226398 7608
rect 277394 7556 277400 7608
rect 277452 7596 277458 7608
rect 332686 7596 332692 7608
rect 277452 7568 332692 7596
rect 277452 7556 277458 7568
rect 332686 7556 332692 7568
rect 332744 7556 332750 7608
rect 335354 7556 335360 7608
rect 335412 7596 335418 7608
rect 481726 7596 481732 7608
rect 335412 7568 481732 7596
rect 335412 7556 335418 7568
rect 481726 7556 481732 7568
rect 481784 7556 481790 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 170398 6848 170404 6860
rect 3476 6820 170404 6848
rect 3476 6808 3482 6820
rect 170398 6808 170404 6820
rect 170456 6808 170462 6860
rect 190362 6808 190368 6860
rect 190420 6848 190426 6860
rect 580166 6848 580172 6860
rect 190420 6820 580172 6848
rect 190420 6808 190426 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 292574 6536 292580 6588
rect 292632 6576 292638 6588
rect 371694 6576 371700 6588
rect 292632 6548 371700 6576
rect 292632 6536 292638 6548
rect 371694 6536 371700 6548
rect 371752 6536 371758 6588
rect 293954 6468 293960 6520
rect 294012 6508 294018 6520
rect 375282 6508 375288 6520
rect 294012 6480 375288 6508
rect 294012 6468 294018 6480
rect 375282 6468 375288 6480
rect 375340 6468 375346 6520
rect 295334 6400 295340 6452
rect 295392 6440 295398 6452
rect 378870 6440 378876 6452
rect 295392 6412 378876 6440
rect 295392 6400 295398 6412
rect 378870 6400 378876 6412
rect 378928 6400 378934 6452
rect 300854 6332 300860 6384
rect 300912 6372 300918 6384
rect 393038 6372 393044 6384
rect 300912 6344 393044 6372
rect 300912 6332 300918 6344
rect 393038 6332 393044 6344
rect 393096 6332 393102 6384
rect 362954 6264 362960 6316
rect 363012 6304 363018 6316
rect 552658 6304 552664 6316
rect 363012 6276 552664 6304
rect 363012 6264 363018 6276
rect 552658 6264 552664 6276
rect 552716 6264 552722 6316
rect 288434 6196 288440 6248
rect 288492 6236 288498 6248
rect 361114 6236 361120 6248
rect 288492 6208 361120 6236
rect 288492 6196 288498 6208
rect 361114 6196 361120 6208
rect 361172 6196 361178 6248
rect 369854 6196 369860 6248
rect 369912 6236 369918 6248
rect 570322 6236 570328 6248
rect 369912 6208 570328 6236
rect 369912 6196 369918 6208
rect 570322 6196 570328 6208
rect 570380 6196 570386 6248
rect 291194 6128 291200 6180
rect 291252 6168 291258 6180
rect 368198 6168 368204 6180
rect 291252 6140 368204 6168
rect 291252 6128 291258 6140
rect 368198 6128 368204 6140
rect 368256 6128 368262 6180
rect 371234 6128 371240 6180
rect 371292 6168 371298 6180
rect 573910 6168 573916 6180
rect 371292 6140 573916 6168
rect 371292 6128 371298 6140
rect 573910 6128 573916 6140
rect 573968 6128 573974 6180
rect 274634 5312 274640 5364
rect 274692 5352 274698 5364
rect 325602 5352 325608 5364
rect 274692 5324 325608 5352
rect 274692 5312 274698 5324
rect 325602 5312 325608 5324
rect 325660 5312 325666 5364
rect 276014 5244 276020 5296
rect 276072 5284 276078 5296
rect 329190 5284 329196 5296
rect 276072 5256 329196 5284
rect 276072 5244 276078 5256
rect 329190 5244 329196 5256
rect 329248 5244 329254 5296
rect 349154 5244 349160 5296
rect 349212 5284 349218 5296
rect 517146 5284 517152 5296
rect 349212 5256 517152 5284
rect 349212 5244 349218 5256
rect 517146 5244 517152 5256
rect 517204 5244 517210 5296
rect 278774 5176 278780 5228
rect 278832 5216 278838 5228
rect 336274 5216 336280 5228
rect 278832 5188 336280 5216
rect 278832 5176 278838 5188
rect 336274 5176 336280 5188
rect 336332 5176 336338 5228
rect 350534 5176 350540 5228
rect 350592 5216 350598 5228
rect 520734 5216 520740 5228
rect 350592 5188 520740 5216
rect 350592 5176 350598 5188
rect 520734 5176 520740 5188
rect 520792 5176 520798 5228
rect 280154 5108 280160 5160
rect 280212 5148 280218 5160
rect 339862 5148 339868 5160
rect 280212 5120 339868 5148
rect 280212 5108 280218 5120
rect 339862 5108 339868 5120
rect 339920 5108 339926 5160
rect 353294 5108 353300 5160
rect 353352 5148 353358 5160
rect 527818 5148 527824 5160
rect 353352 5120 527824 5148
rect 353352 5108 353358 5120
rect 527818 5108 527824 5120
rect 527876 5108 527882 5160
rect 281534 5040 281540 5092
rect 281592 5080 281598 5092
rect 343358 5080 343364 5092
rect 281592 5052 343364 5080
rect 281592 5040 281598 5052
rect 343358 5040 343364 5052
rect 343416 5040 343422 5092
rect 354674 5040 354680 5092
rect 354732 5080 354738 5092
rect 531314 5080 531320 5092
rect 354732 5052 531320 5080
rect 354732 5040 354738 5052
rect 531314 5040 531320 5052
rect 531372 5040 531378 5092
rect 282914 4972 282920 5024
rect 282972 5012 282978 5024
rect 346946 5012 346952 5024
rect 282972 4984 346952 5012
rect 282972 4972 282978 4984
rect 346946 4972 346952 4984
rect 347004 4972 347010 5024
rect 356054 4972 356060 5024
rect 356112 5012 356118 5024
rect 534902 5012 534908 5024
rect 356112 4984 534908 5012
rect 356112 4972 356118 4984
rect 534902 4972 534908 4984
rect 534960 4972 534966 5024
rect 284294 4904 284300 4956
rect 284352 4944 284358 4956
rect 350442 4944 350448 4956
rect 284352 4916 350448 4944
rect 284352 4904 284358 4916
rect 350442 4904 350448 4916
rect 350500 4904 350506 4956
rect 357434 4904 357440 4956
rect 357492 4944 357498 4956
rect 538398 4944 538404 4956
rect 357492 4916 538404 4944
rect 357492 4904 357498 4916
rect 538398 4904 538404 4916
rect 538456 4904 538462 4956
rect 194410 4836 194416 4888
rect 194468 4876 194474 4888
rect 223574 4876 223580 4888
rect 194468 4848 223580 4876
rect 194468 4836 194474 4848
rect 223574 4836 223580 4848
rect 223632 4836 223638 4888
rect 285674 4836 285680 4888
rect 285732 4876 285738 4888
rect 354030 4876 354036 4888
rect 285732 4848 354036 4876
rect 285732 4836 285738 4848
rect 354030 4836 354036 4848
rect 354088 4836 354094 4888
rect 358814 4836 358820 4888
rect 358872 4876 358878 4888
rect 541986 4876 541992 4888
rect 358872 4848 541992 4876
rect 358872 4836 358878 4848
rect 541986 4836 541992 4848
rect 542044 4836 542050 4888
rect 128170 4768 128176 4820
rect 128228 4808 128234 4820
rect 195238 4808 195244 4820
rect 128228 4780 195244 4808
rect 128228 4768 128234 4780
rect 195238 4768 195244 4780
rect 195296 4768 195302 4820
rect 287054 4768 287060 4820
rect 287112 4808 287118 4820
rect 357526 4808 357532 4820
rect 287112 4780 357532 4808
rect 287112 4768 287118 4780
rect 357526 4768 357532 4780
rect 357584 4768 357590 4820
rect 360194 4768 360200 4820
rect 360252 4808 360258 4820
rect 545482 4808 545488 4820
rect 360252 4780 545488 4808
rect 360252 4768 360258 4780
rect 545482 4768 545488 4780
rect 545540 4768 545546 4820
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 508498 4088 508504 4140
rect 508556 4128 508562 4140
rect 510062 4128 510068 4140
rect 508556 4100 510068 4128
rect 508556 4088 508562 4100
rect 510062 4088 510068 4100
rect 510120 4088 510126 4140
rect 576118 4088 576124 4140
rect 576176 4128 576182 4140
rect 577406 4128 577412 4140
rect 576176 4100 577412 4128
rect 576176 4088 576182 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 248414 3952 248420 4004
rect 248472 3992 248478 4004
rect 258258 3992 258264 4004
rect 248472 3964 258264 3992
rect 248472 3952 248478 3964
rect 258258 3952 258264 3964
rect 258316 3952 258322 4004
rect 298094 3952 298100 4004
rect 298152 3992 298158 4004
rect 385954 3992 385960 4004
rect 298152 3964 385960 3992
rect 298152 3952 298158 3964
rect 385954 3952 385960 3964
rect 386012 3952 386018 4004
rect 249794 3884 249800 3936
rect 249852 3924 249858 3936
rect 261754 3924 261760 3936
rect 249852 3896 261760 3924
rect 249852 3884 249858 3896
rect 261754 3884 261760 3896
rect 261812 3884 261818 3936
rect 304994 3884 305000 3936
rect 305052 3924 305058 3936
rect 403618 3924 403624 3936
rect 305052 3896 403624 3924
rect 305052 3884 305058 3896
rect 403618 3884 403624 3896
rect 403676 3884 403682 3936
rect 158898 3816 158904 3868
rect 158956 3856 158962 3868
rect 209774 3856 209780 3868
rect 158956 3828 209780 3856
rect 158956 3816 158962 3828
rect 209774 3816 209780 3828
rect 209832 3816 209838 3868
rect 251174 3816 251180 3868
rect 251232 3856 251238 3868
rect 265342 3856 265348 3868
rect 251232 3828 265348 3856
rect 251232 3816 251238 3828
rect 265342 3816 265348 3828
rect 265400 3816 265406 3868
rect 324314 3816 324320 3868
rect 324372 3856 324378 3868
rect 453298 3856 453304 3868
rect 324372 3828 453304 3856
rect 324372 3816 324378 3828
rect 453298 3816 453304 3828
rect 453356 3816 453362 3868
rect 155402 3748 155408 3800
rect 155460 3788 155466 3800
rect 208394 3788 208400 3800
rect 155460 3760 208400 3788
rect 155460 3748 155466 3760
rect 208394 3748 208400 3760
rect 208452 3748 208458 3800
rect 252554 3748 252560 3800
rect 252612 3788 252618 3800
rect 268838 3788 268844 3800
rect 252612 3760 268844 3788
rect 252612 3748 252618 3760
rect 268838 3748 268844 3760
rect 268896 3748 268902 3800
rect 327074 3748 327080 3800
rect 327132 3788 327138 3800
rect 460382 3788 460388 3800
rect 327132 3760 460388 3788
rect 327132 3748 327138 3760
rect 460382 3748 460388 3760
rect 460440 3748 460446 3800
rect 151814 3680 151820 3732
rect 151872 3720 151878 3732
rect 207014 3720 207020 3732
rect 151872 3692 207020 3720
rect 151872 3680 151878 3692
rect 207014 3680 207020 3692
rect 207072 3680 207078 3732
rect 253934 3680 253940 3732
rect 253992 3720 253998 3732
rect 272426 3720 272432 3732
rect 253992 3692 272432 3720
rect 253992 3680 253998 3692
rect 272426 3680 272432 3692
rect 272484 3680 272490 3732
rect 305638 3680 305644 3732
rect 305696 3720 305702 3732
rect 307938 3720 307944 3732
rect 305696 3692 307944 3720
rect 305696 3680 305702 3692
rect 307938 3680 307944 3692
rect 307996 3680 308002 3732
rect 328454 3680 328460 3732
rect 328512 3720 328518 3732
rect 463970 3720 463976 3732
rect 328512 3692 463976 3720
rect 328512 3680 328518 3692
rect 463970 3680 463976 3692
rect 464028 3680 464034 3732
rect 148318 3612 148324 3664
rect 148376 3652 148382 3664
rect 205634 3652 205640 3664
rect 148376 3624 205640 3652
rect 148376 3612 148382 3624
rect 205634 3612 205640 3624
rect 205692 3612 205698 3664
rect 219250 3612 219256 3664
rect 219308 3652 219314 3664
rect 224218 3652 224224 3664
rect 219308 3624 224224 3652
rect 219308 3612 219314 3624
rect 224218 3612 224224 3624
rect 224276 3612 224282 3664
rect 255314 3612 255320 3664
rect 255372 3652 255378 3664
rect 276014 3652 276020 3664
rect 255372 3624 276020 3652
rect 255372 3612 255378 3624
rect 276014 3612 276020 3624
rect 276072 3612 276078 3664
rect 329834 3612 329840 3664
rect 329892 3652 329898 3664
rect 467466 3652 467472 3664
rect 329892 3624 467472 3652
rect 329892 3612 329898 3624
rect 467466 3612 467472 3624
rect 467524 3612 467530 3664
rect 144730 3544 144736 3596
rect 144788 3584 144794 3596
rect 204254 3584 204260 3596
rect 144788 3556 204260 3584
rect 144788 3544 144794 3556
rect 204254 3544 204260 3556
rect 204312 3544 204318 3596
rect 215662 3544 215668 3596
rect 215720 3584 215726 3596
rect 222838 3584 222844 3596
rect 215720 3556 222844 3584
rect 215720 3544 215726 3556
rect 222838 3544 222844 3556
rect 222896 3544 222902 3596
rect 244274 3544 244280 3596
rect 244332 3584 244338 3596
rect 247586 3584 247592 3596
rect 244332 3556 247592 3584
rect 244332 3544 244338 3556
rect 247586 3544 247592 3556
rect 247644 3544 247650 3596
rect 256694 3544 256700 3596
rect 256752 3584 256758 3596
rect 279510 3584 279516 3596
rect 256752 3556 279516 3584
rect 256752 3544 256758 3556
rect 279510 3544 279516 3556
rect 279568 3544 279574 3596
rect 331214 3544 331220 3596
rect 331272 3584 331278 3596
rect 471054 3584 471060 3596
rect 331272 3556 471060 3584
rect 331272 3544 331278 3556
rect 471054 3544 471060 3556
rect 471112 3544 471118 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 15838 3516 15844 3528
rect 1728 3488 15844 3516
rect 1728 3476 1734 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 202874 3516 202880 3528
rect 141292 3488 202880 3516
rect 141292 3476 141298 3488
rect 202874 3476 202880 3488
rect 202932 3476 202938 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 220078 3516 220084 3528
rect 208636 3488 220084 3516
rect 208636 3476 208642 3488
rect 220078 3476 220084 3488
rect 220136 3476 220142 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 228358 3516 228364 3528
rect 226392 3488 228364 3516
rect 226392 3476 226398 3488
rect 228358 3476 228364 3488
rect 228416 3476 228422 3528
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 237374 3516 237380 3528
rect 229888 3488 237380 3516
rect 229888 3476 229894 3488
rect 237374 3476 237380 3488
rect 237432 3476 237438 3528
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 241514 3516 241520 3528
rect 240560 3488 241520 3516
rect 240560 3476 240566 3488
rect 241514 3476 241520 3488
rect 241572 3476 241578 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244090 3516 244096 3528
rect 242952 3488 244096 3516
rect 242952 3476 242958 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 245654 3476 245660 3528
rect 245712 3516 245718 3528
rect 251174 3516 251180 3528
rect 245712 3488 251180 3516
rect 245712 3476 245718 3488
rect 251174 3476 251180 3488
rect 251232 3476 251238 3528
rect 258074 3476 258080 3528
rect 258132 3516 258138 3528
rect 283098 3516 283104 3528
rect 258132 3488 283104 3516
rect 258132 3476 258138 3488
rect 283098 3476 283104 3488
rect 283156 3476 283162 3528
rect 287698 3476 287704 3528
rect 287756 3516 287762 3528
rect 290182 3516 290188 3528
rect 287756 3488 290188 3516
rect 287756 3476 287762 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 300762 3516 300768 3528
rect 299532 3488 300768 3516
rect 299532 3476 299538 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 309778 3476 309784 3528
rect 309836 3516 309842 3528
rect 311434 3516 311440 3528
rect 309836 3488 311440 3516
rect 309836 3476 309842 3488
rect 311434 3476 311440 3488
rect 311492 3476 311498 3528
rect 333974 3476 333980 3528
rect 334032 3516 334038 3528
rect 478138 3516 478144 3528
rect 334032 3488 478144 3516
rect 334032 3476 334038 3488
rect 478138 3476 478144 3488
rect 478196 3476 478202 3528
rect 494698 3476 494704 3528
rect 494756 3516 494762 3528
rect 495894 3516 495900 3528
rect 494756 3488 495900 3516
rect 494756 3476 494762 3488
rect 495894 3476 495900 3488
rect 495952 3476 495958 3528
rect 512638 3476 512644 3528
rect 512696 3516 512702 3528
rect 513558 3516 513564 3528
rect 512696 3488 513564 3516
rect 512696 3476 512702 3488
rect 513558 3476 513564 3488
rect 513616 3476 513622 3528
rect 555418 3476 555424 3528
rect 555476 3516 555482 3528
rect 556154 3516 556160 3528
rect 555476 3488 556160 3516
rect 555476 3476 555482 3488
rect 556154 3476 556160 3488
rect 556212 3476 556218 3528
rect 137646 3408 137652 3460
rect 137704 3448 137710 3460
rect 201586 3448 201592 3460
rect 137704 3420 201592 3448
rect 137704 3408 137710 3420
rect 201586 3408 201592 3420
rect 201644 3408 201650 3460
rect 205082 3408 205088 3460
rect 205140 3448 205146 3460
rect 218698 3448 218704 3460
rect 205140 3420 218704 3448
rect 205140 3408 205146 3420
rect 218698 3408 218704 3420
rect 218756 3408 218762 3460
rect 222746 3408 222752 3460
rect 222804 3448 222810 3460
rect 233878 3448 233884 3460
rect 222804 3420 233884 3448
rect 222804 3408 222810 3420
rect 233878 3408 233884 3420
rect 233936 3408 233942 3460
rect 247034 3408 247040 3460
rect 247092 3448 247098 3460
rect 254670 3448 254676 3460
rect 247092 3420 254676 3448
rect 247092 3408 247098 3420
rect 254670 3408 254676 3420
rect 254728 3408 254734 3460
rect 259454 3408 259460 3460
rect 259512 3448 259518 3460
rect 286594 3448 286600 3460
rect 259512 3420 286600 3448
rect 259512 3408 259518 3420
rect 286594 3408 286600 3420
rect 286652 3408 286658 3460
rect 373994 3408 374000 3460
rect 374052 3448 374058 3460
rect 580994 3448 581000 3460
rect 374052 3420 581000 3448
rect 374052 3408 374058 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 233418 3204 233424 3256
rect 233476 3244 233482 3256
rect 238754 3244 238760 3256
rect 233476 3216 238760 3244
rect 233476 3204 233482 3216
rect 238754 3204 238760 3216
rect 238812 3204 238818 3256
rect 578878 3204 578884 3256
rect 578936 3244 578942 3256
rect 582190 3244 582196 3256
rect 578936 3216 582196 3244
rect 578936 3204 578942 3216
rect 582190 3204 582196 3216
rect 582248 3204 582254 3256
rect 237006 3000 237012 3052
rect 237064 3040 237070 3052
rect 239398 3040 239404 3052
rect 237064 3012 239404 3040
rect 237064 3000 237070 3012
rect 239398 3000 239404 3012
rect 239456 3000 239462 3052
rect 291930 3000 291936 3052
rect 291988 3040 291994 3052
rect 293678 3040 293684 3052
rect 291988 3012 293684 3040
rect 291988 3000 291994 3012
rect 293678 3000 293684 3012
rect 293736 3000 293742 3052
rect 294046 2864 294052 2916
rect 294104 2904 294110 2916
rect 297266 2904 297272 2916
rect 294104 2876 297272 2904
rect 294104 2864 294110 2876
rect 297266 2864 297272 2876
rect 297324 2864 297330 2916
rect 483658 2864 483664 2916
rect 483716 2904 483722 2916
rect 485222 2904 485228 2916
rect 483716 2876 485228 2904
rect 483716 2864 483722 2876
rect 485222 2864 485228 2876
rect 485280 2864 485286 2916
rect 558178 2864 558184 2916
rect 558236 2904 558242 2916
rect 559742 2904 559748 2916
rect 558236 2876 559748 2904
rect 558236 2864 558242 2876
rect 559742 2864 559748 2876
rect 559800 2864 559806 2916
rect 562318 2864 562324 2916
rect 562376 2904 562382 2916
rect 566826 2904 566832 2916
rect 562376 2876 566832 2904
rect 562376 2864 562382 2876
rect 566826 2864 566832 2876
rect 566884 2864 566890 2916
rect 423674 2728 423680 2780
rect 423732 2768 423738 2780
rect 424962 2768 424968 2780
rect 423732 2740 424968 2768
rect 423732 2728 423738 2740
rect 424962 2728 424968 2740
rect 425020 2728 425026 2780
rect 448514 2728 448520 2780
rect 448572 2768 448578 2780
rect 449802 2768 449808 2780
rect 448572 2740 449808 2768
rect 448572 2728 448578 2740
rect 449802 2728 449808 2740
rect 449860 2728 449866 2780
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 154120 700340 154172 700392
rect 199384 700340 199436 700392
rect 202788 700340 202840 700392
rect 203524 700340 203576 700392
rect 371884 700340 371936 700392
rect 478512 700340 478564 700392
rect 89168 700272 89220 700324
rect 206284 700272 206336 700324
rect 212540 700272 212592 700324
rect 413652 700272 413704 700324
rect 418804 700272 418856 700324
rect 429844 700272 429896 700324
rect 479524 700272 479576 700324
rect 527180 700272 527232 700324
rect 8116 699660 8168 699712
rect 10324 699660 10376 699712
rect 345664 699660 345716 699712
rect 348792 699660 348844 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 558184 699660 558236 699712
rect 559656 699660 559708 699712
rect 215300 697552 215352 697604
rect 218980 697552 219032 697604
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 271144 696940 271196 696992
rect 580172 696940 580224 696992
rect 23480 692044 23532 692096
rect 219440 692044 219492 692096
rect 71780 690616 71832 690668
rect 218060 690616 218112 690668
rect 136640 689256 136692 689308
rect 216680 689256 216732 689308
rect 40040 687896 40092 687948
rect 218152 687896 218204 687948
rect 104900 686468 104952 686520
rect 216772 686468 216824 686520
rect 169760 685108 169812 685160
rect 216864 685108 216916 685160
rect 166448 684904 166500 684956
rect 249800 684904 249852 684956
rect 163964 684836 164016 684888
rect 248420 684836 248472 684888
rect 159272 684768 159324 684820
rect 244280 684768 244332 684820
rect 156880 684700 156932 684752
rect 242900 684700 242952 684752
rect 154304 684632 154356 684684
rect 240140 684632 240192 684684
rect 132960 684564 133012 684616
rect 252560 684564 252612 684616
rect 118608 684496 118660 684548
rect 241520 684496 241572 684548
rect 161388 684020 161440 684072
rect 245660 684020 245712 684072
rect 142160 683952 142212 684004
rect 242992 683952 243044 684004
rect 133880 683884 133932 683936
rect 248512 683884 248564 683936
rect 130384 683816 130436 683868
rect 247040 683816 247092 683868
rect 124220 683748 124272 683800
rect 243084 683748 243136 683800
rect 111064 683680 111116 683732
rect 241612 683680 241664 683732
rect 104256 683612 104308 683664
rect 244372 683612 244424 683664
rect 97080 683544 97132 683596
rect 238760 683544 238812 683596
rect 94688 683476 94740 683528
rect 237656 683476 237708 683528
rect 92296 683408 92348 683460
rect 236000 683408 236052 683460
rect 70768 683340 70820 683392
rect 252652 683340 252704 683392
rect 44180 683272 44232 683324
rect 241704 683272 241756 683324
rect 32496 683204 32548 683256
rect 238852 683204 238904 683256
rect 3424 683136 3476 683188
rect 202144 683136 202196 683188
rect 224224 683136 224276 683188
rect 580172 683136 580224 683188
rect 61200 682864 61252 682916
rect 146944 682864 146996 682916
rect 42064 682796 42116 682848
rect 142160 682796 142212 682848
rect 85120 682728 85172 682780
rect 137284 682728 137336 682780
rect 99288 682660 99340 682712
rect 111064 682660 111116 682712
rect 106648 682592 106700 682644
rect 130384 682592 130436 682644
rect 171048 682592 171100 682644
rect 252744 682592 252796 682644
rect 101864 682524 101916 682576
rect 124220 682524 124272 682576
rect 149704 682524 149756 682576
rect 198188 682524 198240 682576
rect 108948 682456 109000 682508
rect 133880 682456 133932 682508
rect 144828 682456 144880 682508
rect 198280 682456 198332 682508
rect 142528 682388 142580 682440
rect 198004 682388 198056 682440
rect 130568 682320 130620 682372
rect 198096 682320 198148 682372
rect 44088 682252 44140 682304
rect 168380 682252 168432 682304
rect 185584 682252 185636 682304
rect 260840 682252 260892 682304
rect 65984 682184 66036 682236
rect 100760 682184 100812 682236
rect 183192 682184 183244 682236
rect 259736 682184 259788 682236
rect 58808 682116 58860 682168
rect 107568 682116 107620 682168
rect 140136 682116 140188 682168
rect 173808 682116 173860 682168
rect 178408 682116 178460 682168
rect 256700 682116 256752 682168
rect 79968 682048 80020 682100
rect 144276 682048 144328 682100
rect 180616 682048 180668 682100
rect 258356 682048 258408 682100
rect 63408 681980 63460 682032
rect 169760 681980 169812 682032
rect 176016 681980 176068 682032
rect 255320 681980 255372 682032
rect 147312 681912 147364 681964
rect 259552 681912 259604 681964
rect 25320 681844 25372 681896
rect 60740 681844 60792 681896
rect 73068 681844 73120 681896
rect 85488 681844 85540 681896
rect 128176 681844 128228 681896
rect 249892 681844 249944 681896
rect 27528 681776 27580 681828
rect 79048 681776 79100 681828
rect 125416 681776 125468 681828
rect 247224 681776 247276 681828
rect 37188 681708 37240 681760
rect 44180 681708 44232 681760
rect 87512 681708 87564 681760
rect 98644 681708 98696 681760
rect 173624 681708 173676 681760
rect 198372 681708 198424 681760
rect 168380 681300 168432 681352
rect 243176 681300 243228 681352
rect 173808 681232 173860 681284
rect 256792 681232 256844 681284
rect 146944 681164 146996 681216
rect 249984 681164 250036 681216
rect 107568 681096 107620 681148
rect 248696 681096 248748 681148
rect 100760 681028 100812 681080
rect 251180 681028 251232 681080
rect 85488 680960 85540 681012
rect 254216 680960 254268 681012
rect 123392 680824 123444 680876
rect 245844 680824 245896 680876
rect 111432 680756 111484 680808
rect 236184 680756 236236 680808
rect 82728 680688 82780 680740
rect 256884 680688 256936 680740
rect 77944 680620 77996 680672
rect 255412 680620 255464 680672
rect 68376 680552 68428 680604
rect 252836 680552 252888 680604
rect 56416 680484 56468 680536
rect 248604 680484 248656 680536
rect 49240 680416 49292 680468
rect 245752 680416 245804 680468
rect 39672 680348 39724 680400
rect 241796 680348 241848 680400
rect 137284 679668 137336 679720
rect 258172 679668 258224 679720
rect 98644 679600 98696 679652
rect 258264 679600 258316 679652
rect 89720 679396 89772 679448
rect 113824 679396 113876 679448
rect 116032 679396 116084 679448
rect 121000 679396 121052 679448
rect 135168 679396 135220 679448
rect 151912 679396 151964 679448
rect 187792 679396 187844 679448
rect 234712 679396 234764 679448
rect 238944 679328 238996 679380
rect 254032 679260 254084 679312
rect 244556 679192 244608 679244
rect 240324 679124 240376 679176
rect 239036 679056 239088 679108
rect 259644 678988 259696 679040
rect 3516 670692 3568 670744
rect 20904 670692 20956 670744
rect 231124 670692 231176 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 11704 656888 11756 656940
rect 233884 643084 233936 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 208400 630640 208452 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 19984 618264 20036 618316
rect 222844 616836 222896 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 14464 605820 14516 605872
rect 228364 590656 228416 590708
rect 579804 590656 579856 590708
rect 209780 588548 209832 588600
rect 542360 588548 542412 588600
rect 211160 587120 211212 587172
rect 462320 587120 462372 587172
rect 209872 585760 209924 585812
rect 479524 585760 479576 585812
rect 551008 585148 551060 585200
rect 557540 585148 557592 585200
rect 211252 584400 211304 584452
rect 494060 584400 494112 584452
rect 3332 579640 3384 579692
rect 18604 579640 18656 579692
rect 562324 563048 562376 563100
rect 580172 563048 580224 563100
rect 3332 553392 3384 553444
rect 15844 553392 15896 553444
rect 406292 536800 406344 536852
rect 416780 536800 416832 536852
rect 563704 536800 563756 536852
rect 579896 536800 579948 536852
rect 270500 535440 270552 535492
rect 416780 535440 416832 535492
rect 416044 532788 416096 532840
rect 418068 532788 418120 532840
rect 280804 532720 280856 532772
rect 417056 532720 417108 532772
rect 414664 530000 414716 530052
rect 417424 530000 417476 530052
rect 279424 529932 279476 529984
rect 417700 529932 417752 529984
rect 2964 527144 3016 527196
rect 7564 527144 7616 527196
rect 295984 527144 296036 527196
rect 417700 527144 417752 527196
rect 565084 524424 565136 524476
rect 580172 524424 580224 524476
rect 558276 510620 558328 510672
rect 580172 510620 580224 510672
rect 277584 509260 277636 509312
rect 417608 509260 417660 509312
rect 298744 507832 298796 507884
rect 416780 507832 416832 507884
rect 213920 507084 213972 507136
rect 345664 507084 345716 507136
rect 211344 505724 211396 505776
rect 371884 505724 371936 505776
rect 214012 504364 214064 504416
rect 331220 504364 331272 504416
rect 212632 502936 212684 502988
rect 364340 502936 364392 502988
rect 212724 501576 212776 501628
rect 396724 501576 396776 501628
rect 3332 500964 3384 501016
rect 20076 500964 20128 501016
rect 211436 500216 211488 500268
rect 418804 500216 418856 500268
rect 205640 498788 205692 498840
rect 558276 498788 558328 498840
rect 551928 498176 551980 498228
rect 557540 498176 557592 498228
rect 476764 498040 476816 498092
rect 480352 498040 480404 498092
rect 65248 497428 65300 497480
rect 151084 497428 151136 497480
rect 276020 497224 276072 497276
rect 485780 497224 485832 497276
rect 283564 497156 283616 497208
rect 452660 497156 452712 497208
rect 262220 497088 262272 497140
rect 436192 497088 436244 497140
rect 260932 497020 260984 497072
rect 436100 497020 436152 497072
rect 457444 497020 457496 497072
rect 473360 497020 473412 497072
rect 277492 496952 277544 497004
rect 459560 496952 459612 497004
rect 464344 496952 464396 497004
rect 476120 496952 476172 497004
rect 271880 496884 271932 496936
rect 470784 496884 470836 496936
rect 475384 496884 475436 496936
rect 483020 496884 483072 496936
rect 472624 496816 472676 496868
rect 477500 496816 477552 496868
rect 269120 496136 269172 496188
rect 448520 496136 448572 496188
rect 274640 496068 274692 496120
rect 455420 496068 455472 496120
rect 262312 494708 262364 494760
rect 437480 494708 437532 494760
rect 273260 493280 273312 493332
rect 454040 493280 454092 493332
rect 215392 491988 215444 492040
rect 282920 491988 282972 492040
rect 276112 491920 276164 491972
rect 458272 491920 458324 491972
rect 274732 490560 274784 490612
rect 456892 490560 456944 490612
rect 276204 489200 276256 489252
rect 456800 489200 456852 489252
rect 205732 489132 205784 489184
rect 562324 489132 562376 489184
rect 262404 487772 262456 487824
rect 443092 487772 443144 487824
rect 266452 486412 266504 486464
rect 441620 486412 441672 486464
rect 226984 484372 227036 484424
rect 580172 484372 580224 484424
rect 263600 483624 263652 483676
rect 438860 483624 438912 483676
rect 209964 482332 210016 482384
rect 224224 482332 224276 482384
rect 3516 482264 3568 482316
rect 223580 482264 223632 482316
rect 271972 482264 272024 482316
rect 467840 482264 467892 482316
rect 3424 480972 3476 481024
rect 222200 480972 222252 481024
rect 270592 480972 270644 481024
rect 465080 480972 465132 481024
rect 207020 480904 207072 480956
rect 580264 480904 580316 480956
rect 19984 479544 20036 479596
rect 220820 479544 220872 479596
rect 269212 479544 269264 479596
rect 460940 479544 460992 479596
rect 205824 479476 205876 479528
rect 565084 479476 565136 479528
rect 208492 478184 208544 478236
rect 271144 478184 271196 478236
rect 21364 478116 21416 478168
rect 220912 478116 220964 478168
rect 269304 478116 269356 478168
rect 462320 478116 462372 478168
rect 206284 476892 206336 476944
rect 218244 476892 218296 476944
rect 214104 476824 214156 476876
rect 266360 476824 266412 476876
rect 22100 476756 22152 476808
rect 236276 476756 236328 476808
rect 267740 476756 267792 476808
rect 458180 476756 458232 476808
rect 266360 475328 266412 475380
rect 454684 475328 454736 475380
rect 3424 474716 3476 474768
rect 223672 474716 223724 474768
rect 20076 474036 20128 474088
rect 223764 474036 223816 474088
rect 264980 474036 265032 474088
rect 452752 474036 452804 474088
rect 205916 473968 205968 474020
rect 563704 473968 563756 474020
rect 214196 472676 214248 472728
rect 299480 472676 299532 472728
rect 15844 472608 15896 472660
rect 222292 472608 222344 472660
rect 263692 472608 263744 472660
rect 449992 472608 450044 472660
rect 14464 471248 14516 471300
rect 221004 471248 221056 471300
rect 270684 471248 270736 471300
rect 451372 471248 451424 471300
rect 204260 470568 204312 470620
rect 579988 470568 580040 470620
rect 207112 469888 207164 469940
rect 228364 469888 228416 469940
rect 270776 469888 270828 469940
rect 449900 469888 449952 469940
rect 11704 469820 11756 469872
rect 219532 469820 219584 469872
rect 273352 469820 273404 469872
rect 464344 469820 464396 469872
rect 204352 468528 204404 468580
rect 226984 468528 227036 468580
rect 267832 468528 267884 468580
rect 447232 468528 447284 468580
rect 10324 468460 10376 468512
rect 219624 468460 219676 468512
rect 273444 468460 273496 468512
rect 457444 468460 457496 468512
rect 208584 467168 208636 467220
rect 233884 467168 233936 467220
rect 261024 467168 261076 467220
rect 298744 467168 298796 467220
rect 7564 467100 7616 467152
rect 222384 467100 222436 467152
rect 276296 467100 276348 467152
rect 475384 467100 475436 467152
rect 198924 466828 198976 466880
rect 577688 466828 577740 466880
rect 198832 466760 198884 466812
rect 577872 466760 577924 466812
rect 198740 466692 198792 466744
rect 577964 466692 578016 466744
rect 200120 466624 200172 466676
rect 580540 466624 580592 466676
rect 197636 466556 197688 466608
rect 577780 466556 577832 466608
rect 196072 466488 196124 466540
rect 577504 466488 577556 466540
rect 196164 466420 196216 466472
rect 580264 466420 580316 466472
rect 269396 465808 269448 465860
rect 280804 465808 280856 465860
rect 18604 465740 18656 465792
rect 222476 465740 222528 465792
rect 274824 465740 274876 465792
rect 472624 465740 472676 465792
rect 210056 465672 210108 465724
rect 558184 465672 558236 465724
rect 160744 465468 160796 465520
rect 367100 465468 367152 465520
rect 161020 465400 161072 465452
rect 370136 465400 370188 465452
rect 160928 465332 160980 465384
rect 372620 465332 372672 465384
rect 160836 465264 160888 465316
rect 375380 465264 375432 465316
rect 14648 465196 14700 465248
rect 231952 465196 232004 465248
rect 197452 465128 197504 465180
rect 577596 465128 577648 465180
rect 197544 465060 197596 465112
rect 580356 465060 580408 465112
rect 169024 464584 169076 464636
rect 327356 464584 327408 464636
rect 316316 464516 316368 464568
rect 395344 464516 395396 464568
rect 199384 464448 199436 464500
rect 216956 464448 217008 464500
rect 302240 464448 302292 464500
rect 394056 464448 394108 464500
rect 208676 464380 208728 464432
rect 231124 464380 231176 464432
rect 267924 464380 267976 464432
rect 416044 464380 416096 464432
rect 4804 464312 4856 464364
rect 221096 464312 221148 464364
rect 266544 464312 266596 464364
rect 445760 464312 445812 464364
rect 320364 464244 320416 464296
rect 406200 464244 406252 464296
rect 166724 464176 166776 464228
rect 331496 464176 331548 464228
rect 166356 464108 166408 464160
rect 333980 464108 334032 464160
rect 166816 464040 166868 464092
rect 336740 464040 336792 464092
rect 166540 463972 166592 464024
rect 341156 463972 341208 464024
rect 166448 463904 166500 463956
rect 343640 463904 343692 463956
rect 166264 463836 166316 463888
rect 346584 463836 346636 463888
rect 171784 463768 171836 463820
rect 380900 463768 380952 463820
rect 199016 463700 199068 463752
rect 580448 463700 580500 463752
rect 174636 463292 174688 463344
rect 378140 463292 378192 463344
rect 202144 463224 202196 463276
rect 219716 463224 219768 463276
rect 266636 463224 266688 463276
rect 279424 463224 279476 463276
rect 159732 463156 159784 463208
rect 294144 463156 294196 463208
rect 349252 463156 349304 463208
rect 407856 463156 407908 463208
rect 159640 463088 159692 463140
rect 298192 463088 298244 463140
rect 346492 463088 346544 463140
rect 410616 463088 410668 463140
rect 159364 463020 159416 463072
rect 302332 463020 302384 463072
rect 342260 463020 342312 463072
rect 410708 463020 410760 463072
rect 167736 462952 167788 463004
rect 233516 462952 233568 463004
rect 261116 462952 261168 463004
rect 447140 462952 447192 463004
rect 159548 462884 159600 462936
rect 306380 462884 306432 462936
rect 336832 462884 336884 462936
rect 407764 462884 407816 462936
rect 309140 462816 309192 462868
rect 395436 462816 395488 462868
rect 159456 462748 159508 462800
rect 314660 462748 314712 462800
rect 330116 462748 330168 462800
rect 408040 462748 408092 462800
rect 162124 462680 162176 462732
rect 317420 462680 317472 462732
rect 323124 462680 323176 462732
rect 405004 462680 405056 462732
rect 161112 462612 161164 462664
rect 310520 462612 310572 462664
rect 339500 462612 339552 462664
rect 407948 462612 408000 462664
rect 174544 462544 174596 462596
rect 375472 462544 375524 462596
rect 163688 462476 163740 462528
rect 351920 462476 351972 462528
rect 354772 462476 354824 462528
rect 410800 462476 410852 462528
rect 14556 462408 14608 462460
rect 232044 462408 232096 462460
rect 305000 462408 305052 462460
rect 403624 462408 403676 462460
rect 3240 462340 3292 462392
rect 225144 462340 225196 462392
rect 298284 462340 298336 462392
rect 416044 462340 416096 462392
rect 177304 461932 177356 461984
rect 342352 461932 342404 461984
rect 167920 461864 167972 461916
rect 229100 461864 229152 461916
rect 195980 461796 196032 461848
rect 196164 461796 196216 461848
rect 203524 461796 203576 461848
rect 215576 461796 215628 461848
rect 161204 461728 161256 461780
rect 290004 461728 290056 461780
rect 313280 461728 313332 461780
rect 395528 461728 395580 461780
rect 207204 461660 207256 461712
rect 222844 461660 222896 461712
rect 265072 461660 265124 461712
rect 414664 461660 414716 461712
rect 215484 461592 215536 461644
rect 234620 461592 234672 461644
rect 245660 461592 245712 461644
rect 246396 461592 246448 461644
rect 263784 461592 263836 461644
rect 443000 461592 443052 461644
rect 334072 461524 334124 461576
rect 400772 461524 400824 461576
rect 177488 461456 177540 461508
rect 347780 461456 347832 461508
rect 174820 461388 174872 461440
rect 357440 461388 357492 461440
rect 174912 461320 174964 461372
rect 362960 461320 363012 461372
rect 174728 461252 174780 461304
rect 368480 461252 368532 461304
rect 204444 461184 204496 461236
rect 559564 461184 559616 461236
rect 202880 461116 202932 461168
rect 558276 461116 558328 461168
rect 201500 461048 201552 461100
rect 563704 461048 563756 461100
rect 202972 460980 203024 461032
rect 576124 460980 576176 461032
rect 203064 460912 203116 460964
rect 580724 460912 580776 460964
rect 237564 460776 237616 460828
rect 237932 460776 237984 460828
rect 177396 460572 177448 460624
rect 354864 460572 354916 460624
rect 169300 460504 169352 460556
rect 280988 460504 281040 460556
rect 167828 460436 167880 460488
rect 231308 460436 231360 460488
rect 264428 460436 264480 460488
rect 295984 460436 296036 460488
rect 316132 460436 316184 460488
rect 405372 460436 405424 460488
rect 172060 460368 172112 460420
rect 297548 460368 297600 460420
rect 318800 460368 318852 460420
rect 411812 460368 411864 460420
rect 171968 460300 172020 460352
rect 301596 460300 301648 460352
rect 309232 460300 309284 460352
rect 405280 460300 405332 460352
rect 198372 460232 198424 460284
rect 254492 460232 254544 460284
rect 272156 460232 272208 460284
rect 451280 460232 451332 460284
rect 275468 460164 275520 460216
rect 476764 460164 476816 460216
rect 301044 460096 301096 460148
rect 402520 460096 402572 460148
rect 177672 460028 177724 460080
rect 345756 460028 345808 460080
rect 356796 460028 356848 460080
rect 400956 460028 401008 460080
rect 164148 459960 164200 460012
rect 338396 459960 338448 460012
rect 396724 459960 396776 460012
rect 171876 459892 171928 459944
rect 305644 459892 305696 459944
rect 350908 459892 350960 459944
rect 401048 459892 401100 459944
rect 14924 459824 14976 459876
rect 230572 459824 230624 459876
rect 292764 459824 292816 459876
rect 402244 459824 402296 459876
rect 14464 459756 14516 459808
rect 233332 459756 233384 459808
rect 286508 459756 286560 459808
rect 418896 459756 418948 459808
rect 159824 459688 159876 459740
rect 385500 459688 385552 459740
rect 156696 459620 156748 459672
rect 382556 459620 382608 459672
rect 204536 459552 204588 459604
rect 493416 459552 493468 459604
rect 240140 459484 240192 459536
rect 240876 459484 240928 459536
rect 185676 459280 185728 459332
rect 336188 459280 336240 459332
rect 188528 459212 188580 459264
rect 319628 459212 319680 459264
rect 162492 459144 162544 459196
rect 328552 459144 328604 459196
rect 198188 459076 198240 459128
rect 237380 459076 237432 459128
rect 283656 459076 283708 459128
rect 400864 459076 400916 459128
rect 198096 459008 198148 459060
rect 251364 459008 251416 459060
rect 353852 459008 353904 459060
rect 401140 459008 401192 459060
rect 198004 458940 198056 458992
rect 258080 458940 258132 458992
rect 347964 458940 348016 458992
rect 401232 458940 401284 458992
rect 188896 458872 188948 458924
rect 299664 458872 299716 458924
rect 305184 458872 305236 458924
rect 402428 458872 402480 458924
rect 197360 458804 197412 458856
rect 197544 458804 197596 458856
rect 198280 458804 198332 458856
rect 259460 458804 259512 458856
rect 265532 458804 265584 458856
rect 444380 458804 444432 458856
rect 252836 458736 252888 458788
rect 253020 458736 253072 458788
rect 287980 458736 288032 458788
rect 402336 458736 402388 458788
rect 221004 458668 221056 458720
rect 221372 458668 221424 458720
rect 296812 458668 296864 458720
rect 402612 458668 402664 458720
rect 216772 458600 216824 458652
rect 217692 458600 217744 458652
rect 219532 458600 219584 458652
rect 220268 458600 220320 458652
rect 312636 458600 312688 458652
rect 405464 458600 405516 458652
rect 188620 458532 188672 458584
rect 323124 458532 323176 458584
rect 325700 458532 325752 458584
rect 403992 458532 404044 458584
rect 188344 458464 188396 458516
rect 329932 458464 329984 458516
rect 332692 458464 332744 458516
rect 415308 458464 415360 458516
rect 186964 458396 187016 458448
rect 291200 458396 291252 458448
rect 329196 458396 329248 458448
rect 403900 458396 403952 458448
rect 177580 458328 177632 458380
rect 339868 458328 339920 458380
rect 342444 458328 342496 458380
rect 404084 458328 404136 458380
rect 187056 458260 187108 458312
rect 303988 458260 304040 458312
rect 319260 458260 319312 458312
rect 418804 458260 418856 458312
rect 15016 458192 15068 458244
rect 230664 458192 230716 458244
rect 369952 458192 370004 458244
rect 413376 458192 413428 458244
rect 493416 458124 493468 458176
rect 580172 458124 580224 458176
rect 180616 457852 180668 457904
rect 326620 457852 326672 457904
rect 162400 457784 162452 457836
rect 361948 457784 362000 457836
rect 162768 457716 162820 457768
rect 359004 457716 359056 457768
rect 180432 457648 180484 457700
rect 333244 457648 333296 457700
rect 356428 457648 356480 457700
rect 412364 457648 412416 457700
rect 183284 457580 183336 457632
rect 288440 457580 288492 457632
rect 289268 457580 289320 457632
rect 354220 457580 354272 457632
rect 372712 457580 372764 457632
rect 416136 457580 416188 457632
rect 180340 457512 180392 457564
rect 292856 457512 292908 457564
rect 359372 457512 359424 457564
rect 411996 457512 412048 457564
rect 170496 457444 170548 457496
rect 234988 457444 235040 457496
rect 265256 457444 265308 457496
rect 440240 457444 440292 457496
rect 180248 457376 180300 457428
rect 297180 457376 297232 457428
rect 338764 457376 338816 457428
rect 412456 457376 412508 457428
rect 180156 457308 180208 457360
rect 301228 457308 301280 457360
rect 335452 457308 335504 457360
rect 412272 457308 412324 457360
rect 318984 457240 319036 457292
rect 414664 457240 414716 457292
rect 278688 457172 278740 457224
rect 419264 457172 419316 457224
rect 325976 457104 326028 457156
rect 414756 457104 414808 457156
rect 308588 457036 308640 457088
rect 406568 457036 406620 457088
rect 180524 456968 180576 457020
rect 320180 456968 320232 457020
rect 332140 456968 332192 457020
rect 414848 456968 414900 457020
rect 169392 456900 169444 456952
rect 316684 456900 316736 456952
rect 341708 456900 341760 456952
rect 412088 456900 412140 456952
rect 172152 456832 172204 456884
rect 288716 456832 288768 456884
rect 348056 456832 348108 456884
rect 412180 456832 412232 456884
rect 162308 456764 162360 456816
rect 364892 456764 364944 456816
rect 375288 456764 375340 456816
rect 388904 456764 388956 456816
rect 162676 456560 162728 456612
rect 370780 456560 370832 456612
rect 216680 456492 216732 456544
rect 216956 456492 217008 456544
rect 219440 456492 219492 456544
rect 219716 456492 219768 456544
rect 244280 456492 244332 456544
rect 244648 456492 244700 456544
rect 328552 456492 328604 456544
rect 414572 456492 414624 456544
rect 165160 456424 165212 456476
rect 374092 456424 374144 456476
rect 162584 456356 162636 456408
rect 367836 456356 367888 456408
rect 172244 456288 172296 456340
rect 293408 456288 293460 456340
rect 333980 456288 334032 456340
rect 334348 456288 334400 456340
rect 377036 456288 377088 456340
rect 409328 456288 409380 456340
rect 167644 456220 167696 456272
rect 234252 456220 234304 456272
rect 276020 456220 276072 456272
rect 276940 456220 276992 456272
rect 282184 456220 282236 456272
rect 416320 456220 416372 456272
rect 188804 456152 188856 456204
rect 279516 456152 279568 456204
rect 282460 456152 282512 456204
rect 419356 456152 419408 456204
rect 200764 456084 200816 456136
rect 331220 456084 331272 456136
rect 336740 456084 336792 456136
rect 337660 456084 337712 456136
rect 354680 456084 354732 456136
rect 355692 456084 355744 456136
rect 375380 456084 375432 456136
rect 376300 456084 376352 456136
rect 376392 456084 376444 456136
rect 398104 456084 398156 456136
rect 165068 456016 165120 456068
rect 311440 456016 311492 456068
rect 352380 456016 352432 456068
rect 395620 456016 395672 456068
rect 215300 455948 215352 456000
rect 216220 455948 216272 456000
rect 218152 455948 218204 456000
rect 218796 455948 218848 456000
rect 220820 455948 220872 456000
rect 221740 455948 221792 456000
rect 222384 455948 222436 456000
rect 223212 455948 223264 456000
rect 223672 455948 223724 456000
rect 224316 455948 224368 456000
rect 231952 455948 232004 456000
rect 232780 455948 232832 456000
rect 244372 455948 244424 456000
rect 244924 455948 244976 456000
rect 247224 455948 247276 456000
rect 247868 455948 247920 456000
rect 251180 455948 251232 456000
rect 251916 455948 251968 456000
rect 252652 455948 252704 456000
rect 253388 455948 253440 456000
rect 273352 455948 273404 456000
rect 273996 455948 274048 456000
rect 276112 455948 276164 456000
rect 276572 455948 276624 456000
rect 312268 455948 312320 456000
rect 403716 455948 403768 456000
rect 164056 455880 164108 455932
rect 316316 455880 316368 455932
rect 339132 455880 339184 455932
rect 404176 455880 404228 455932
rect 191196 455812 191248 455864
rect 200764 455812 200816 455864
rect 322204 455812 322256 455864
rect 414940 455812 414992 455864
rect 158076 455744 158128 455796
rect 330024 455744 330076 455796
rect 374460 455744 374512 455796
rect 376392 455744 376444 455796
rect 158260 455676 158312 455728
rect 322940 455676 322992 455728
rect 358268 455676 358320 455728
rect 392952 455676 393004 455728
rect 273444 455608 273496 455660
rect 273628 455608 273680 455660
rect 368664 455608 368716 455660
rect 409236 455608 409288 455660
rect 162216 455540 162268 455592
rect 313372 455540 313424 455592
rect 371516 455540 371568 455592
rect 398196 455540 398248 455592
rect 164976 455472 165028 455524
rect 376760 455472 376812 455524
rect 377404 455472 377456 455524
rect 398288 455472 398340 455524
rect 164884 455404 164936 455456
rect 379888 455404 379940 455456
rect 381728 455404 381780 455456
rect 416228 455404 416280 455456
rect 18972 455064 19024 455116
rect 299480 455064 299532 455116
rect 19064 454996 19116 455048
rect 295984 454996 296036 455048
rect 306656 454996 306708 455048
rect 394332 454996 394384 455048
rect 188988 454928 189040 454980
rect 278044 454928 278096 454980
rect 278688 454928 278740 454980
rect 328828 454928 328880 454980
rect 415032 454928 415084 454980
rect 166908 454860 166960 454912
rect 285956 454860 286008 454912
rect 317512 454860 317564 454912
rect 388536 454860 388588 454912
rect 191288 454792 191340 454844
rect 321836 454792 321888 454844
rect 169484 454724 169536 454776
rect 309968 454724 310020 454776
rect 331220 454792 331272 454844
rect 331772 454792 331824 454844
rect 389916 454792 389968 454844
rect 396816 454724 396868 454776
rect 168104 454656 168156 454708
rect 310520 454656 310572 454708
rect 314108 454656 314160 454708
rect 394148 454656 394200 454708
rect 172336 454588 172388 454640
rect 344560 454588 344612 454640
rect 169668 454520 169720 454572
rect 347504 454520 347556 454572
rect 363144 454520 363196 454572
rect 401324 454520 401376 454572
rect 161296 454452 161348 454504
rect 353300 454452 353352 454504
rect 361212 454452 361264 454504
rect 418988 454452 419040 454504
rect 14832 454384 14884 454436
rect 230940 454384 230992 454436
rect 285036 454384 285088 454436
rect 391296 454384 391348 454436
rect 289452 454316 289504 454368
rect 391388 454316 391440 454368
rect 294144 454248 294196 454300
rect 391204 454248 391256 454300
rect 18880 454180 18932 454232
rect 304080 454180 304132 454232
rect 304724 454180 304776 454232
rect 310704 454180 310756 454232
rect 394240 454180 394292 454232
rect 18788 454112 18840 454164
rect 308128 454112 308180 454164
rect 375932 454112 375984 454164
rect 392768 454112 392820 454164
rect 19340 454044 19392 454096
rect 312176 454044 312228 454096
rect 384304 454044 384356 454096
rect 389364 454044 389416 454096
rect 175096 453636 175148 453688
rect 341616 453636 341668 453688
rect 347872 453636 347924 453688
rect 348056 453636 348108 453688
rect 17408 453568 17460 453620
rect 291660 453568 291712 453620
rect 304724 453568 304776 453620
rect 417516 453568 417568 453620
rect 214104 453500 214156 453552
rect 214748 453500 214800 453552
rect 258264 453500 258316 453552
rect 258908 453500 258960 453552
rect 269304 453500 269356 453552
rect 269948 453500 270000 453552
rect 273168 453500 273220 453552
rect 283564 453500 283616 453552
rect 299480 453500 299532 453552
rect 300032 453500 300084 453552
rect 390284 453500 390336 453552
rect 191472 453432 191524 453484
rect 282460 453432 282512 453484
rect 295984 453432 296036 453484
rect 390192 453432 390244 453484
rect 189816 453364 189868 453416
rect 325056 453364 325108 453416
rect 343824 453364 343876 453416
rect 182732 453296 182784 453348
rect 328368 453296 328420 453348
rect 340880 453296 340932 453348
rect 179972 453228 180024 453280
rect 331680 453228 331732 453280
rect 177212 453160 177264 453212
rect 338120 453160 338172 453212
rect 342260 453160 342312 453212
rect 343180 453160 343232 453212
rect 349160 453160 349212 453212
rect 349804 453160 349856 453212
rect 371240 453296 371292 453348
rect 375288 453296 375340 453348
rect 395804 453228 395856 453280
rect 395896 453160 395948 453212
rect 191380 453092 191432 453144
rect 356060 453092 356112 453144
rect 364340 453092 364392 453144
rect 393136 453092 393188 453144
rect 17776 453024 17828 453076
rect 4068 452956 4120 453008
rect 226064 452956 226116 453008
rect 234712 452956 234764 453008
rect 235356 452956 235408 453008
rect 236092 452956 236144 453008
rect 236552 452956 236604 453008
rect 237472 452956 237524 453008
rect 238300 452956 238352 453008
rect 238944 452956 238996 453008
rect 239128 452956 239180 453008
rect 241520 452956 241572 453008
rect 242348 452956 242400 453008
rect 242992 452956 243044 453008
rect 243452 452956 243504 453008
rect 254124 452956 254176 453008
rect 254860 452956 254912 453008
rect 255320 452956 255372 453008
rect 255964 452956 256016 453008
rect 256792 452956 256844 453008
rect 257068 452956 257120 453008
rect 258080 452956 258132 453008
rect 258264 452956 258316 453008
rect 259552 452956 259604 453008
rect 260380 452956 260432 453008
rect 260932 452956 260984 453008
rect 261484 452956 261536 453008
rect 262220 452956 262272 453008
rect 262956 452956 263008 453008
rect 263600 452956 263652 453008
rect 263784 452956 263836 453008
rect 269120 452956 269172 453008
rect 269304 452956 269356 453008
rect 270684 452956 270736 453008
rect 271420 452956 271472 453008
rect 271880 452956 271932 453008
rect 272524 452956 272576 453008
rect 3424 452888 3476 452940
rect 227536 452888 227588 452940
rect 236184 452888 236236 452940
rect 236828 452888 236880 452940
rect 238760 452888 238812 452940
rect 239404 452888 239456 452940
rect 256700 452888 256752 452940
rect 257436 452888 257488 452940
rect 259644 452888 259696 452940
rect 260012 452888 260064 452940
rect 270592 452888 270644 452940
rect 271052 452888 271104 452940
rect 302332 453024 302384 453076
rect 302700 453024 302752 453076
rect 337568 453024 337620 453076
rect 398656 453024 398708 453076
rect 291660 452956 291712 453008
rect 390100 452956 390152 453008
rect 287152 452888 287204 452940
rect 388812 452888 388864 452940
rect 3332 452820 3384 452872
rect 226432 452820 226484 452872
rect 238852 452820 238904 452872
rect 239772 452820 239824 452872
rect 312176 452820 312228 452872
rect 417700 452820 417752 452872
rect 3792 452752 3844 452804
rect 228640 452752 228692 452804
rect 308128 452752 308180 452804
rect 417608 452752 417660 452804
rect 198740 452684 198792 452736
rect 199292 452684 199344 452736
rect 202880 452684 202932 452736
rect 203708 452684 203760 452736
rect 204352 452684 204404 452736
rect 204812 452684 204864 452736
rect 205824 452684 205876 452736
rect 206284 452684 206336 452736
rect 207020 452684 207072 452736
rect 207388 452684 207440 452736
rect 208492 452684 208544 452736
rect 209228 452684 209280 452736
rect 209872 452684 209924 452736
rect 210332 452684 210384 452736
rect 211160 452684 211212 452736
rect 211436 452684 211488 452736
rect 212540 452684 212592 452736
rect 212908 452684 212960 452736
rect 213920 452684 213972 452736
rect 214104 452684 214156 452736
rect 287520 452684 287572 452736
rect 416964 452684 417016 452736
rect 193864 452616 193916 452668
rect 224960 452616 225012 452668
rect 370320 452616 370372 452668
rect 392860 452616 392912 452668
rect 198832 452548 198884 452600
rect 199660 452548 199712 452600
rect 204260 452548 204312 452600
rect 205180 452548 205232 452600
rect 205732 452548 205784 452600
rect 206652 452548 206704 452600
rect 209780 452548 209832 452600
rect 210700 452548 210752 452600
rect 212632 452548 212684 452600
rect 213276 452548 213328 452600
rect 299664 452480 299716 452532
rect 303896 452480 303948 452532
rect 156972 452208 157024 452260
rect 294880 452208 294932 452260
rect 163412 452140 163464 452192
rect 303712 452140 303764 452192
rect 304264 452140 304316 452192
rect 367376 452276 367428 452328
rect 375196 452276 375248 452328
rect 385040 452276 385092 452328
rect 394424 452276 394476 452328
rect 325424 452208 325476 452260
rect 387708 452208 387760 452260
rect 335360 452140 335412 452192
rect 336648 452140 336700 452192
rect 349712 452140 349764 452192
rect 371240 452140 371292 452192
rect 378784 452140 378836 452192
rect 385224 452140 385276 452192
rect 188252 452072 188304 452124
rect 286508 452072 286560 452124
rect 291200 452072 291252 452124
rect 297364 452072 297416 452124
rect 303988 452072 304040 452124
rect 397184 452072 397236 452124
rect 191012 452004 191064 452056
rect 290464 452004 290516 452056
rect 303896 452004 303948 452056
rect 397092 452004 397144 452056
rect 189908 451936 189960 451988
rect 295616 451936 295668 451988
rect 297640 451936 297692 451988
rect 190000 451868 190052 451920
rect 297824 451868 297876 451920
rect 303712 451868 303764 451920
rect 304264 451936 304316 451988
rect 396908 451936 396960 451988
rect 307760 451868 307812 451920
rect 397000 451868 397052 451920
rect 191748 451800 191800 451852
rect 314752 451800 314804 451852
rect 320824 451800 320876 451852
rect 378784 451800 378836 451852
rect 380992 451800 381044 451852
rect 381176 451800 381228 451852
rect 157800 451732 157852 451784
rect 282368 451732 282420 451784
rect 297364 451732 297416 451784
rect 394516 451732 394568 451784
rect 158628 451664 158680 451716
rect 286416 451664 286468 451716
rect 413836 451664 413888 451716
rect 190920 451596 190972 451648
rect 318800 451596 318852 451648
rect 336648 451596 336700 451648
rect 388720 451596 388772 451648
rect 208308 451528 208360 451580
rect 208584 451528 208636 451580
rect 253940 451528 253992 451580
rect 254216 451528 254268 451580
rect 282368 451528 282420 451580
rect 413744 451528 413796 451580
rect 158352 451460 158404 451512
rect 282184 451460 282236 451512
rect 290832 451460 290884 451512
rect 416504 451460 416556 451512
rect 156880 451392 156932 451444
rect 299296 451392 299348 451444
rect 314752 451392 314804 451444
rect 315488 451392 315540 451444
rect 320824 451392 320876 451444
rect 158444 451324 158496 451376
rect 325424 451324 325476 451376
rect 187608 451256 187660 451308
rect 196992 451256 197044 451308
rect 210516 451256 210568 451308
rect 222476 451256 222528 451308
rect 222660 451256 222712 451308
rect 225696 451256 225748 451308
rect 278780 451256 278832 451308
rect 296352 451256 296404 451308
rect 310520 451256 310572 451308
rect 311808 451256 311860 451308
rect 417424 451392 417476 451444
rect 375196 451324 375248 451376
rect 393044 451324 393096 451376
rect 373264 451256 373316 451308
rect 419080 451256 419132 451308
rect 166172 451052 166224 451104
rect 350448 451052 350500 451104
rect 279424 450984 279476 451036
rect 389824 450984 389876 451036
rect 280896 450916 280948 450968
rect 409696 450916 409748 450968
rect 210424 450848 210476 450900
rect 375104 450848 375156 450900
rect 191656 450780 191708 450832
rect 281632 450780 281684 450832
rect 177948 450712 178000 450764
rect 284576 450712 284628 450764
rect 298192 450712 298244 450764
rect 298652 450712 298704 450764
rect 168196 450644 168248 450696
rect 295248 450644 295300 450696
rect 298560 450644 298612 450696
rect 394608 450712 394660 450764
rect 368848 450644 368900 450696
rect 398564 450644 398616 450696
rect 3240 450576 3292 450628
rect 210516 450576 210568 450628
rect 320640 450576 320692 450628
rect 382188 450576 382240 450628
rect 17868 450508 17920 450560
rect 278780 450508 278832 450560
rect 293776 450508 293828 450560
rect 358728 450508 358780 450560
rect 365904 450508 365956 450560
rect 401416 450508 401468 450560
rect 186136 450440 186188 450492
rect 321744 450440 321796 450492
rect 365536 450440 365588 450492
rect 409512 450440 409564 450492
rect 191564 450372 191616 450424
rect 334992 450372 335044 450424
rect 336096 450372 336148 450424
rect 403532 450372 403584 450424
rect 186044 450304 186096 450356
rect 339776 450304 339828 450356
rect 346768 450304 346820 450356
rect 395712 450304 395764 450356
rect 191840 450236 191892 450288
rect 222108 450236 222160 450288
rect 222200 450236 222252 450288
rect 222844 450236 222896 450288
rect 223580 450236 223632 450288
rect 223948 450236 224000 450288
rect 244464 450236 244516 450288
rect 245292 450236 245344 450288
rect 249800 450236 249852 450288
rect 250076 450236 250128 450288
rect 252560 450236 252612 450288
rect 252928 450236 252980 450288
rect 274732 450236 274784 450288
rect 275100 450236 275152 450288
rect 302240 450236 302292 450288
rect 302424 450236 302476 450288
rect 322940 450236 322992 450288
rect 323308 450236 323360 450288
rect 362960 450236 363012 450288
rect 363420 450236 363472 450288
rect 371424 450236 371476 450288
rect 409420 450236 409472 450288
rect 177856 450168 177908 450220
rect 351920 450168 351972 450220
rect 362592 450168 362644 450220
rect 412548 450168 412600 450220
rect 222292 450100 222344 450152
rect 227168 450100 227220 450152
rect 345296 450100 345348 450152
rect 404268 450100 404320 450152
rect 165252 450032 165304 450084
rect 290556 450032 290608 450084
rect 383476 450032 383528 450084
rect 407028 450032 407080 450084
rect 3976 449964 4028 450016
rect 226616 449964 226668 450016
rect 270500 449964 270552 450016
rect 270776 449964 270828 450016
rect 325700 449964 325752 450016
rect 325976 449964 326028 450016
rect 374276 449964 374328 450016
rect 409604 449964 409656 450016
rect 19248 449896 19300 449948
rect 278504 449896 278556 449948
rect 380808 449896 380860 449948
rect 398472 449896 398524 449948
rect 190828 449828 190880 449880
rect 193864 449828 193916 449880
rect 193956 449828 194008 449880
rect 201224 449828 201276 449880
rect 3700 449692 3752 449744
rect 200856 449692 200908 449744
rect 382280 449760 382332 449812
rect 3884 449624 3936 449676
rect 193128 449624 193180 449676
rect 193220 449624 193272 449676
rect 195336 449624 195388 449676
rect 228088 449692 228140 449744
rect 382740 449692 382792 449744
rect 386420 449692 386472 449744
rect 386512 449692 386564 449744
rect 387616 449692 387668 449744
rect 387708 449692 387760 449744
rect 388996 449692 389048 449744
rect 413928 449692 413980 449744
rect 165344 449556 165396 449608
rect 3516 449488 3568 449540
rect 190828 449488 190880 449540
rect 200856 449556 200908 449608
rect 201224 449556 201276 449608
rect 379428 449624 379480 449676
rect 416688 449624 416740 449676
rect 307208 449556 307260 449608
rect 336740 449556 336792 449608
rect 385224 449556 385276 449608
rect 385684 449556 385736 449608
rect 388076 449556 388128 449608
rect 399484 449556 399536 449608
rect 388996 449488 389048 449540
rect 411076 449488 411128 449540
rect 131764 444728 131816 444780
rect 134340 444728 134392 444780
rect 151084 435344 151136 435396
rect 158720 435344 158772 435396
rect 551928 435344 551980 435396
rect 557540 435344 557592 435396
rect 19156 433984 19208 434036
rect 131764 433984 131816 434036
rect 154580 433984 154632 434036
rect 184204 433984 184256 434036
rect 558276 431876 558328 431928
rect 580080 431876 580132 431928
rect 559564 419432 559616 419484
rect 580080 419432 580132 419484
rect 563796 405628 563848 405680
rect 580080 405628 580132 405680
rect 388904 384956 388956 385008
rect 390376 384956 390428 385008
rect 17500 384276 17552 384328
rect 18880 384276 18932 384328
rect 390284 382916 390336 382968
rect 416780 382916 416832 382968
rect 17684 382236 17736 382288
rect 18972 382236 19024 382288
rect 390192 381488 390244 381540
rect 416872 381488 416924 381540
rect 390100 380128 390152 380180
rect 416780 380128 416832 380180
rect 576124 379448 576176 379500
rect 580080 379448 580132 379500
rect 388904 378768 388956 378820
rect 416780 378768 416832 378820
rect 558184 353200 558236 353252
rect 580080 353200 580132 353252
rect 399484 349868 399536 349920
rect 418160 349868 418212 349920
rect 390376 349800 390428 349852
rect 492588 349800 492640 349852
rect 103520 349596 103572 349648
rect 162768 349596 162820 349648
rect 418160 349596 418212 349648
rect 419448 349596 419500 349648
rect 452568 349596 452620 349648
rect 98552 349528 98604 349580
rect 161296 349528 161348 349580
rect 408224 349528 408276 349580
rect 478512 349528 478564 349580
rect 93492 349460 93544 349512
rect 169668 349460 169720 349512
rect 400772 349460 400824 349512
rect 483480 349460 483532 349512
rect 91008 349392 91060 349444
rect 172336 349392 172388 349444
rect 398656 349392 398708 349444
rect 485964 349392 486016 349444
rect 78036 349324 78088 349376
rect 163412 349324 163464 349376
rect 395896 349324 395948 349376
rect 488264 349324 488316 349376
rect 71780 349256 71832 349308
rect 72240 349256 72292 349308
rect 190920 349256 190972 349308
rect 395804 349256 395856 349308
rect 491024 349256 491076 349308
rect 67640 349188 67692 349240
rect 68744 349188 68796 349240
rect 190000 349188 190052 349240
rect 416688 349188 416740 349240
rect 520924 349188 520976 349240
rect 62856 349120 62908 349172
rect 188252 349120 188304 349172
rect 393136 349120 393188 349172
rect 508504 349120 508556 349172
rect 62028 349052 62080 349104
rect 157800 349052 157852 349104
rect 388904 349052 388956 349104
rect 419540 349052 419592 349104
rect 61108 348984 61160 349036
rect 158536 348984 158588 349036
rect 414572 348984 414624 349036
rect 418068 348984 418120 349036
rect 58532 348916 58584 348968
rect 156880 348916 156932 348968
rect 56048 348848 56100 348900
rect 156972 348848 157024 348900
rect 78496 348780 78548 348832
rect 182732 348780 182784 348832
rect 420000 348780 420052 348832
rect 500960 348780 501012 348832
rect 50804 348712 50856 348764
rect 166908 348712 166960 348764
rect 418988 348712 419040 348764
rect 505928 348712 505980 348764
rect 39580 348644 39632 348696
rect 158628 348644 158680 348696
rect 411076 348644 411128 348696
rect 418712 348644 418764 348696
rect 419080 348644 419132 348696
rect 515864 348644 515916 348696
rect 38476 348576 38528 348628
rect 158352 348576 158404 348628
rect 395620 348576 395672 348628
rect 498476 348576 498528 348628
rect 71136 348508 71188 348560
rect 190828 348508 190880 348560
rect 413928 348508 413980 348560
rect 523316 348508 523368 348560
rect 65156 348440 65208 348492
rect 189908 348440 189960 348492
rect 392952 348440 393004 348492
rect 503444 348440 503496 348492
rect 53656 348372 53708 348424
rect 190920 348372 190972 348424
rect 393044 348372 393096 348424
rect 510988 348372 511040 348424
rect 86040 348304 86092 348356
rect 177212 348304 177264 348356
rect 68376 348236 68428 348288
rect 157892 348236 157944 348288
rect 73160 348168 73212 348220
rect 74356 348168 74408 348220
rect 158444 348168 158496 348220
rect 418712 347896 418764 347948
rect 455788 347896 455840 347948
rect 19156 347828 19208 347880
rect 38476 347828 38528 347880
rect 419540 347828 419592 347880
rect 458180 347828 458232 347880
rect 18696 347760 18748 347812
rect 39580 347760 39632 347812
rect 418068 347760 418120 347812
rect 456984 347760 457036 347812
rect 462228 347760 462280 347812
rect 42800 347692 42852 347744
rect 62028 347692 62080 347744
rect 64788 347692 64840 347744
rect 186964 347692 187016 347744
rect 417424 347692 417476 347744
rect 417976 347692 418028 347744
rect 458180 347692 458232 347744
rect 459468 347692 459520 347744
rect 478052 347692 478104 347744
rect 45928 347624 45980 347676
rect 46572 347624 46624 347676
rect 65156 347624 65208 347676
rect 66260 347624 66312 347676
rect 188896 347624 188948 347676
rect 394608 347624 394660 347676
rect 458364 347624 458416 347676
rect 462228 347624 462280 347676
rect 475660 347624 475712 347676
rect 477408 347624 477460 347676
rect 479156 347624 479208 347676
rect 44180 347556 44232 347608
rect 62856 347556 62908 347608
rect 67732 347556 67784 347608
rect 187056 347556 187108 347608
rect 391388 347556 391440 347608
rect 453580 347556 453632 347608
rect 455788 347556 455840 347608
rect 474372 347556 474424 347608
rect 51080 347488 51132 347540
rect 52368 347488 52420 347540
rect 71136 347488 71188 347540
rect 73252 347488 73304 347540
rect 190828 347488 190880 347540
rect 391296 347488 391348 347540
rect 450636 347488 450688 347540
rect 452568 347488 452620 347540
rect 471244 347488 471296 347540
rect 16488 347216 16540 347268
rect 53472 347420 53524 347472
rect 71780 347420 71832 347472
rect 76748 347420 76800 347472
rect 190920 347420 190972 347472
rect 409696 347420 409748 347472
rect 448244 347420 448296 347472
rect 50068 347352 50120 347404
rect 67640 347352 67692 347404
rect 76104 347352 76156 347404
rect 189816 347352 189868 347404
rect 416320 347352 416372 347404
rect 418896 347352 418948 347404
rect 419356 347352 419408 347404
rect 437020 347352 437072 347404
rect 73712 347284 73764 347336
rect 186136 347284 186188 347336
rect 411812 347284 411864 347336
rect 419724 347284 419776 347336
rect 436744 347284 436796 347336
rect 443092 347284 443144 347336
rect 461492 347284 461544 347336
rect 56600 347216 56652 347268
rect 73160 347216 73212 347268
rect 83648 347216 83700 347268
rect 190828 347216 190880 347268
rect 413836 347216 413888 347268
rect 419172 347216 419224 347268
rect 419264 347216 419316 347268
rect 436100 347216 436152 347268
rect 452568 347216 452620 347268
rect 469772 347216 469824 347268
rect 45376 347148 45428 347200
rect 19616 347080 19668 347132
rect 37188 347080 37240 347132
rect 19892 347012 19944 347064
rect 42800 347012 42852 347064
rect 19800 346944 19852 346996
rect 44180 346944 44232 346996
rect 18972 346876 19024 346928
rect 64788 347148 64840 347200
rect 81072 347148 81124 347200
rect 179972 347148 180024 347200
rect 419080 347148 419132 347200
rect 49608 347080 49660 347132
rect 67732 347080 67784 347132
rect 100944 347080 100996 347132
rect 190920 347080 190972 347132
rect 389916 347080 389968 347132
rect 419632 347080 419684 347132
rect 419816 347080 419868 347132
rect 440516 347080 440568 347132
rect 456800 347148 456852 347200
rect 458088 347148 458140 347200
rect 476948 347148 477000 347200
rect 444196 347080 444248 347132
rect 462780 347080 462832 347132
rect 18604 346808 18656 346860
rect 45928 346808 45980 346860
rect 16120 346740 16172 346792
rect 47584 346740 47636 346792
rect 66260 347012 66312 347064
rect 75460 347012 75512 347064
rect 162492 347012 162544 347064
rect 417976 347012 418028 347064
rect 451372 347012 451424 347064
rect 452568 347012 452620 347064
rect 453028 347012 453080 347064
rect 472072 347012 472124 347064
rect 60832 346944 60884 346996
rect 78036 346944 78088 346996
rect 79140 346944 79192 346996
rect 164148 346944 164200 346996
rect 391204 346944 391256 346996
rect 456156 346944 456208 346996
rect 125968 346876 126020 346928
rect 159824 346876 159876 346928
rect 416504 346876 416556 346928
rect 419816 346876 419868 346928
rect 123392 346808 123444 346860
rect 156696 346808 156748 346860
rect 419632 346808 419684 346860
rect 456800 346808 456852 346860
rect 448520 346740 448572 346792
rect 467380 346740 467432 346792
rect 18236 346672 18288 346724
rect 16212 346604 16264 346656
rect 48596 346604 48648 346656
rect 49608 346604 49660 346656
rect 16304 346536 16356 346588
rect 50068 346536 50120 346588
rect 55220 346672 55272 346724
rect 73252 346672 73304 346724
rect 447140 346672 447192 346724
rect 465724 346672 465776 346724
rect 59360 346604 59412 346656
rect 76748 346604 76800 346656
rect 446404 346604 446456 346656
rect 465172 346604 465224 346656
rect 51264 346536 51316 346588
rect 69296 346536 69348 346588
rect 419172 346536 419224 346588
rect 439596 346536 439648 346588
rect 445300 346536 445352 346588
rect 463884 346536 463936 346588
rect 16396 346468 16448 346520
rect 51080 346468 51132 346520
rect 61936 346468 61988 346520
rect 79140 346468 79192 346520
rect 419724 346468 419776 346520
rect 453028 346468 453080 346520
rect 455236 346468 455288 346520
rect 473360 346468 473412 346520
rect 19708 346400 19760 346452
rect 418896 346400 418948 346452
rect 438032 346400 438084 346452
rect 438860 346400 438912 346452
rect 441620 346400 441672 346452
rect 449900 346400 449952 346452
rect 468668 346400 468720 346452
rect 36176 346332 36228 346384
rect 188988 346332 189040 346384
rect 394424 346332 394476 346384
rect 525892 346332 525944 346384
rect 63684 346264 63736 346316
rect 165344 346264 165396 346316
rect 392768 346264 392820 346316
rect 518348 346264 518400 346316
rect 65984 346196 66036 346248
rect 165068 346196 165120 346248
rect 392860 346196 392912 346248
rect 513380 346196 513432 346248
rect 96068 346128 96120 346180
rect 166172 346128 166224 346180
rect 394240 346128 394292 346180
rect 465264 346128 465316 346180
rect 106096 346060 106148 346112
rect 162400 346060 162452 346112
rect 413744 346060 413796 346112
rect 420000 346060 420052 346112
rect 459560 346060 459612 346112
rect 460572 346060 460624 346112
rect 477408 346060 477460 346112
rect 108672 345992 108724 346044
rect 162308 345992 162360 346044
rect 394056 345992 394108 346044
rect 460940 345992 460992 346044
rect 111064 345924 111116 345976
rect 162584 345924 162636 345976
rect 396908 345924 396960 345976
rect 414572 345924 414624 345976
rect 446404 345924 446456 345976
rect 115848 345856 115900 345908
rect 165160 345856 165212 345908
rect 397184 345856 397236 345908
rect 415860 345856 415912 345908
rect 448520 345856 448572 345908
rect 113456 345788 113508 345840
rect 162676 345788 162728 345840
rect 394516 345788 394568 345840
rect 415952 345788 416004 345840
rect 416688 345788 416740 345840
rect 449900 345788 449952 345840
rect 118608 345720 118660 345772
rect 164976 345720 165028 345772
rect 396816 345720 396868 345772
rect 419908 345720 419960 345772
rect 455236 345720 455288 345772
rect 121000 345652 121052 345704
rect 164884 345652 164936 345704
rect 396724 345652 396776 345704
rect 414480 345652 414532 345704
rect 459560 345652 459612 345704
rect 397092 345584 397144 345636
rect 416320 345584 416372 345636
rect 447140 345584 447192 345636
rect 415952 345516 416004 345568
rect 445300 345516 445352 345568
rect 397000 345448 397052 345500
rect 416688 345448 416740 345500
rect 420000 345448 420052 345500
rect 436744 345448 436796 345500
rect 394332 345312 394384 345364
rect 463516 345312 463568 345364
rect 19984 345040 20036 345092
rect 41328 345040 41380 345092
rect 42708 344972 42760 345024
rect 168196 344972 168248 345024
rect 394148 344972 394200 345024
rect 467932 344972 467984 345024
rect 165252 344904 165304 344956
rect 69296 344836 69348 344888
rect 168104 344836 168156 344888
rect 3424 344292 3476 344344
rect 168012 344292 168064 344344
rect 418620 342932 418672 342984
rect 418896 342932 418948 342984
rect 415860 340144 415912 340196
rect 416504 340144 416556 340196
rect 551008 335452 551060 335504
rect 557540 335452 557592 335504
rect 150992 335316 151044 335368
rect 158720 335248 158772 335300
rect 18880 334908 18932 334960
rect 55220 334908 55272 334960
rect 18328 334840 18380 334892
rect 56600 334840 56652 334892
rect 18788 334772 18840 334824
rect 57980 334772 58032 334824
rect 18512 334704 18564 334756
rect 59360 334704 59412 334756
rect 19524 334636 19576 334688
rect 60740 334636 60792 334688
rect 16028 334568 16080 334620
rect 60832 334568 60884 334620
rect 563704 325592 563756 325644
rect 579620 325592 579672 325644
rect 17040 259360 17092 259412
rect 17316 259360 17368 259412
rect 392676 259360 392728 259412
rect 417884 259360 417936 259412
rect 389916 258068 389968 258120
rect 417148 258068 417200 258120
rect 418620 258068 418672 258120
rect 417700 253172 417752 253224
rect 418620 253172 418672 253224
rect 388168 251812 388220 251864
rect 406292 251812 406344 251864
rect 19340 249704 19392 249756
rect 19616 249704 19668 249756
rect 111064 249704 111116 249756
rect 174452 249704 174504 249756
rect 378232 249704 378284 249756
rect 378784 249704 378836 249756
rect 389916 249704 389968 249756
rect 403532 249704 403584 249756
rect 485964 249704 486016 249756
rect 108580 249636 108632 249688
rect 174912 249636 174964 249688
rect 404176 249636 404228 249688
rect 488264 249636 488316 249688
rect 19432 249568 19484 249620
rect 19708 249568 19760 249620
rect 106004 249568 106056 249620
rect 175188 249568 175240 249620
rect 404084 249568 404136 249620
rect 491024 249568 491076 249620
rect 103520 249500 103572 249552
rect 174820 249500 174872 249552
rect 401232 249500 401284 249552
rect 495900 249500 495952 249552
rect 98552 249432 98604 249484
rect 177856 249432 177908 249484
rect 401048 249432 401100 249484
rect 498476 249432 498528 249484
rect 95884 249364 95936 249416
rect 177488 249364 177540 249416
rect 308588 249364 308640 249416
rect 311164 249364 311216 249416
rect 401140 249364 401192 249416
rect 500960 249364 501012 249416
rect 93492 249296 93544 249348
rect 177672 249296 177724 249348
rect 400956 249296 401008 249348
rect 503536 249296 503588 249348
rect 58532 249228 58584 249280
rect 172060 249228 172112 249280
rect 401508 249228 401560 249280
rect 505928 249228 505980 249280
rect 56048 249160 56100 249212
rect 172244 249160 172296 249212
rect 401324 249160 401376 249212
rect 508504 249160 508556 249212
rect 53656 249092 53708 249144
rect 172152 249092 172204 249144
rect 398196 249092 398248 249144
rect 515864 249092 515916 249144
rect 15752 249024 15804 249076
rect 18604 249024 18656 249076
rect 45928 249024 45980 249076
rect 50804 249024 50856 249076
rect 177948 249024 178000 249076
rect 398288 249024 398340 249076
rect 520924 249024 520976 249076
rect 113456 248956 113508 249008
rect 174728 248956 174780 249008
rect 415308 248956 415360 249008
rect 483480 248956 483532 249008
rect 115848 248888 115900 248940
rect 175004 248888 175056 248940
rect 405372 248888 405424 248940
rect 470968 248888 471020 248940
rect 120908 248820 120960 248872
rect 174636 248820 174688 248872
rect 418804 248820 418856 248872
rect 473636 248820 473688 248872
rect 16304 248344 16356 248396
rect 19708 248412 19760 248464
rect 50160 248344 50212 248396
rect 61200 248344 61252 248396
rect 171968 248344 172020 248396
rect 184204 248344 184256 248396
rect 379612 248344 379664 248396
rect 382372 248344 382424 248396
rect 19248 248276 19300 248328
rect 36452 248276 36504 248328
rect 63592 248276 63644 248328
rect 171876 248276 171928 248328
rect 18604 248208 18656 248260
rect 19432 248208 19484 248260
rect 29552 248208 29604 248260
rect 38660 248208 38712 248260
rect 45928 248208 45980 248260
rect 46664 248208 46716 248260
rect 64880 248208 64932 248260
rect 73804 248208 73856 248260
rect 180524 248208 180576 248260
rect 385132 248344 385184 248396
rect 390652 248344 390704 248396
rect 402244 248276 402296 248328
rect 455420 248276 455472 248328
rect 390560 248208 390612 248260
rect 402336 248208 402388 248260
rect 452660 248208 452712 248260
rect 35900 248140 35952 248192
rect 44180 248140 44232 248192
rect 62120 248140 62172 248192
rect 65984 248140 66036 248192
rect 169484 248140 169536 248192
rect 383752 248140 383804 248192
rect 390744 248140 390796 248192
rect 400864 248140 400916 248192
rect 450360 248140 450412 248192
rect 19156 248072 19208 248124
rect 37280 248072 37332 248124
rect 38108 248072 38160 248124
rect 41420 248072 41472 248124
rect 59452 248072 59504 248124
rect 77300 248072 77352 248124
rect 78496 248072 78548 248124
rect 180616 248072 180668 248124
rect 380992 248072 381044 248124
rect 389180 248072 389232 248124
rect 389824 248072 389876 248124
rect 447140 248072 447192 248124
rect 450176 248072 450228 248124
rect 451280 248072 451332 248124
rect 467840 248072 467892 248124
rect 19984 248004 20036 248056
rect 40040 248004 40092 248056
rect 61384 248004 61436 248056
rect 68376 248004 68428 248056
rect 169576 248004 169628 248056
rect 444472 248004 444524 248056
rect 462320 248004 462372 248056
rect 19892 247936 19944 247988
rect 43076 247936 43128 247988
rect 44272 247936 44324 247988
rect 45284 247936 45336 247988
rect 63500 247936 63552 247988
rect 70952 247936 71004 247988
rect 169392 247936 169444 247988
rect 443184 247936 443236 247988
rect 444196 247936 444248 247988
rect 461124 247936 461176 247988
rect 19800 247868 19852 247920
rect 44180 247868 44232 247920
rect 50160 247868 50212 247920
rect 67640 247868 67692 247920
rect 83648 247868 83700 247920
rect 180432 247868 180484 247920
rect 224224 247868 224276 247920
rect 233332 247868 233384 247920
rect 447140 247868 447192 247920
rect 465080 247868 465132 247920
rect 16120 247800 16172 247852
rect 47584 247800 47636 247852
rect 66260 247800 66312 247852
rect 86040 247800 86092 247852
rect 177764 247800 177816 247852
rect 220084 247800 220136 247852
rect 229192 247800 229244 247852
rect 306472 247800 306524 247852
rect 407120 247800 407172 247852
rect 451372 247800 451424 247852
rect 452476 247800 452528 247852
rect 469220 247800 469272 247852
rect 16212 247732 16264 247784
rect 48688 247732 48740 247784
rect 67732 247732 67784 247784
rect 88248 247732 88300 247784
rect 177580 247732 177632 247784
rect 222844 247732 222896 247784
rect 231952 247732 232004 247784
rect 307852 247732 307904 247784
rect 409880 247732 409932 247784
rect 18512 247664 18564 247716
rect 58072 247664 58124 247716
rect 75920 247664 75972 247716
rect 91008 247664 91060 247716
rect 177304 247664 177356 247716
rect 218704 247664 218756 247716
rect 227812 247664 227864 247716
rect 228364 247664 228416 247716
rect 236092 247664 236144 247716
rect 309232 247664 309284 247716
rect 414020 247664 414072 247716
rect 418528 247664 418580 247716
rect 455880 247732 455932 247784
rect 473360 247732 473412 247784
rect 462228 247664 462280 247716
rect 478880 247664 478932 247716
rect 15660 247596 15712 247648
rect 18972 247596 19024 247648
rect 44272 247596 44324 247648
rect 63224 247596 63276 247648
rect 75000 247596 75052 247648
rect 76104 247596 76156 247648
rect 158260 247596 158312 247648
rect 449900 247596 449952 247648
rect 466460 247596 466512 247648
rect 81072 247528 81124 247580
rect 158076 247528 158128 247580
rect 448520 247528 448572 247580
rect 465080 247528 465132 247580
rect 101220 247460 101272 247512
rect 177396 247460 177448 247512
rect 452752 247460 452804 247512
rect 470784 247460 470836 247512
rect 16028 247392 16080 247444
rect 17040 247392 17092 247444
rect 59452 247392 59504 247444
rect 458272 247392 458324 247444
rect 476120 247392 476172 247444
rect 52552 247324 52604 247376
rect 69020 247324 69072 247376
rect 445760 247324 445812 247376
rect 463700 247324 463752 247376
rect 52460 247256 52512 247308
rect 70400 247256 70452 247308
rect 459560 247256 459612 247308
rect 477500 247256 477552 247308
rect 53840 247188 53892 247240
rect 71780 247188 71832 247240
rect 455420 247188 455472 247240
rect 473360 247188 473412 247240
rect 18512 247120 18564 247172
rect 19340 247120 19392 247172
rect 55128 247120 55180 247172
rect 73160 247120 73212 247172
rect 454040 247120 454092 247172
rect 471980 247120 472032 247172
rect 15936 247052 15988 247104
rect 16212 247052 16264 247104
rect 19064 247052 19116 247104
rect 19248 247052 19300 247104
rect 19432 247052 19484 247104
rect 19984 247052 20036 247104
rect 56600 247052 56652 247104
rect 73252 247052 73304 247104
rect 195244 247052 195296 247104
rect 196072 247052 196124 247104
rect 199384 247052 199436 247104
rect 200212 247052 200264 247104
rect 239404 247052 239456 247104
rect 240232 247052 240284 247104
rect 271972 247052 272024 247104
rect 273904 247052 273956 247104
rect 289912 247052 289964 247104
rect 298744 247052 298796 247104
rect 299572 247052 299624 247104
rect 302884 247052 302936 247104
rect 311992 247052 312044 247104
rect 313924 247052 313976 247104
rect 325792 247052 325844 247104
rect 329104 247052 329156 247104
rect 332692 247052 332744 247104
rect 336004 247052 336056 247104
rect 398380 246984 398432 247036
rect 525800 246984 525852 247036
rect 398564 246916 398616 246968
rect 513380 246916 513432 246968
rect 401416 246848 401468 246900
rect 510620 246848 510672 246900
rect 365812 246372 365864 246424
rect 558184 246372 558236 246424
rect 372712 246304 372764 246356
rect 576124 246304 576176 246356
rect 387064 245624 387116 245676
rect 387892 245624 387944 245676
rect 398472 245556 398524 245608
rect 523040 245556 523092 245608
rect 404268 245488 404320 245540
rect 492680 245488 492732 245540
rect 403900 245420 403952 245472
rect 480536 245420 480588 245472
rect 165620 244944 165672 244996
rect 212632 244944 212684 244996
rect 7564 244876 7616 244928
rect 191932 244876 191984 244928
rect 418620 243516 418672 243568
rect 418988 243516 419040 243568
rect 186320 242156 186372 242208
rect 220912 242156 220964 242208
rect 3516 241408 3568 241460
rect 167920 241408 167972 241460
rect 179420 240728 179472 240780
rect 218060 240728 218112 240780
rect 387064 240728 387116 240780
rect 557632 240728 557684 240780
rect 558828 240728 558880 240780
rect 419632 238688 419684 238740
rect 458272 238688 458324 238740
rect 419816 238620 419868 238672
rect 454040 238620 454092 238672
rect 368480 238076 368532 238128
rect 562324 238076 562376 238128
rect 190184 238008 190236 238060
rect 580540 238008 580592 238060
rect 415860 237396 415912 237448
rect 419632 237396 419684 237448
rect 376760 236648 376812 236700
rect 582380 236648 582432 236700
rect 17316 235900 17368 235952
rect 150440 235900 150492 235952
rect 156696 235900 156748 235952
rect 158628 235900 158680 235952
rect 378784 235900 378836 235952
rect 417700 235900 417752 235952
rect 550824 235900 550876 235952
rect 557448 235900 557500 235952
rect 18328 235832 18380 235884
rect 56600 235832 56652 235884
rect 418068 235832 418120 235884
rect 458180 235832 458232 235884
rect 16304 235764 16356 235816
rect 16488 235764 16540 235816
rect 53840 235764 53892 235816
rect 419908 235764 419960 235816
rect 455420 235764 455472 235816
rect 16028 235696 16080 235748
rect 16396 235696 16448 235748
rect 52460 235696 52512 235748
rect 416688 235696 416740 235748
rect 451280 235696 451332 235748
rect 18880 235628 18932 235680
rect 55220 235628 55272 235680
rect 416504 235628 416556 235680
rect 449900 235628 449952 235680
rect 18236 235560 18288 235612
rect 52552 235560 52604 235612
rect 419448 235560 419500 235612
rect 452752 235560 452804 235612
rect 416320 235492 416372 235544
rect 448520 235492 448572 235544
rect 419080 235424 419132 235476
rect 444472 235424 444524 235476
rect 414572 235356 414624 235408
rect 418988 235356 419040 235408
rect 447140 235356 447192 235408
rect 415952 235288 416004 235340
rect 417148 235288 417200 235340
rect 445760 235288 445812 235340
rect 19524 235220 19576 235272
rect 57980 235220 58032 235272
rect 311164 235220 311216 235272
rect 340144 235220 340196 235272
rect 417976 235220 418028 235272
rect 419540 235220 419592 235272
rect 452660 235220 452712 235272
rect 419724 235152 419776 235204
rect 420000 235152 420052 235204
rect 444380 235152 444432 235204
rect 18236 235084 18288 235136
rect 18696 235084 18748 235136
rect 418712 235084 418764 235136
rect 419356 235084 419408 235136
rect 436100 235084 436152 235136
rect 418896 235016 418948 235068
rect 419264 235016 419316 235068
rect 436192 235016 436244 235068
rect 18788 234948 18840 235000
rect 19524 234948 19576 235000
rect 415676 234744 415728 234796
rect 416504 234744 416556 234796
rect 415768 234676 415820 234728
rect 416688 234676 416740 234728
rect 150440 234608 150492 234660
rect 156696 234608 156748 234660
rect 416320 234608 416372 234660
rect 416504 234608 416556 234660
rect 418436 234608 418488 234660
rect 419080 234608 419132 234660
rect 556804 234540 556856 234592
rect 557540 234540 557592 234592
rect 15844 233860 15896 233912
rect 193220 233860 193272 233912
rect 197360 233860 197412 233912
rect 224960 233860 225012 233912
rect 375380 233860 375432 233912
rect 578884 233860 578936 233912
rect 577964 233180 578016 233232
rect 579620 233180 579672 233232
rect 158720 230392 158772 230444
rect 387064 230392 387116 230444
rect 172520 228352 172572 228404
rect 215300 228352 215352 228404
rect 176660 226992 176712 227044
rect 216680 226992 216732 227044
rect 303620 226992 303672 227044
rect 398840 226992 398892 227044
rect 183560 225564 183612 225616
rect 219440 225564 219492 225616
rect 340144 221076 340196 221128
rect 345112 221076 345164 221128
rect 577872 219172 577924 219224
rect 579988 219172 580040 219224
rect 3332 215228 3384 215280
rect 15108 215228 15160 215280
rect 345112 214548 345164 214600
rect 359464 214548 359516 214600
rect 359464 207612 359516 207664
rect 374644 207612 374696 207664
rect 273904 206252 273956 206304
rect 317512 206252 317564 206304
rect 3056 202784 3108 202836
rect 15016 202784 15068 202836
rect 577780 193128 577832 193180
rect 579620 193128 579672 193180
rect 3516 188980 3568 189032
rect 14924 188980 14976 189032
rect 264980 180072 265032 180124
rect 299480 180072 299532 180124
rect 302240 180072 302292 180124
rect 396080 180072 396132 180124
rect 577688 179324 577740 179376
rect 580080 179324 580132 179376
rect 260840 175924 260892 175976
rect 287704 175924 287756 175976
rect 296720 175924 296772 175976
rect 382280 175924 382332 175976
rect 374644 170280 374696 170332
rect 377220 170280 377272 170332
rect 377220 167968 377272 168020
rect 379520 167968 379572 168020
rect 379520 164840 379572 164892
rect 400864 164840 400916 164892
rect 3240 164160 3292 164212
rect 14832 164160 14884 164212
rect 415216 158108 415268 158160
rect 417700 158108 417752 158160
rect 400864 157972 400916 158024
rect 410984 157972 411036 158024
rect 415860 149676 415912 149728
rect 417700 149676 417752 149728
rect 458088 149676 458140 149728
rect 414756 149608 414808 149660
rect 478512 149608 478564 149660
rect 415032 149540 415084 149592
rect 480904 149540 480956 149592
rect 414848 149472 414900 149524
rect 483480 149472 483532 149524
rect 412272 149404 412324 149456
rect 485964 149404 486016 149456
rect 412456 149336 412508 149388
rect 488264 149336 488316 149388
rect 412088 149268 412140 149320
rect 491024 149268 491076 149320
rect 412180 149200 412232 149252
rect 495900 149200 495952 149252
rect 412364 149132 412416 149184
rect 503536 149132 503588 149184
rect 15108 149064 15160 149116
rect 19616 149064 19668 149116
rect 409604 149064 409656 149116
rect 518440 149064 518492 149116
rect 98552 148996 98604 149048
rect 183468 148996 183520 149048
rect 403716 148996 403768 149048
rect 468300 148996 468352 149048
rect 93492 148928 93544 148980
rect 185952 148928 186004 148980
rect 403808 148928 403860 148980
rect 470968 148928 471020 148980
rect 86040 148860 86092 148912
rect 185676 148860 185728 148912
rect 411996 148860 412048 148912
rect 505928 148860 505980 148912
rect 83556 148792 83608 148844
rect 188712 148792 188764 148844
rect 412548 148792 412600 148844
rect 508504 148792 508556 148844
rect 76104 148724 76156 148776
rect 188620 148724 188672 148776
rect 409512 148724 409564 148776
rect 510988 148724 511040 148776
rect 19616 148656 19668 148708
rect 60648 148656 60700 148708
rect 73620 148656 73672 148708
rect 188528 148656 188580 148708
rect 409236 148656 409288 148708
rect 513380 148656 513432 148708
rect 58532 148588 58584 148640
rect 180248 148588 180300 148640
rect 409420 148588 409472 148640
rect 515864 148588 515916 148640
rect 56048 148520 56100 148572
rect 180340 148520 180392 148572
rect 409328 148520 409380 148572
rect 520924 148520 520976 148572
rect 53656 148452 53708 148504
rect 183284 148452 183336 148504
rect 406936 148452 406988 148504
rect 523316 148452 523368 148504
rect 19708 148384 19760 148436
rect 19984 148384 20036 148436
rect 50804 148384 50856 148436
rect 185860 148384 185912 148436
rect 407028 148384 407080 148436
rect 525892 148384 525944 148436
rect 48320 148316 48372 148368
rect 188804 148316 188856 148368
rect 410984 148316 411036 148368
rect 531044 148316 531096 148368
rect 113456 148248 113508 148300
rect 183100 148248 183152 148300
rect 406568 148248 406620 148300
rect 466000 148248 466052 148300
rect 115848 148180 115900 148232
rect 183008 148180 183060 148232
rect 406752 148180 406804 148232
rect 463516 148180 463568 148232
rect 120908 148112 120960 148164
rect 182824 148112 182876 148164
rect 17040 147840 17092 147892
rect 19708 147840 19760 147892
rect 19984 147840 20036 147892
rect 48228 147840 48280 147892
rect 48136 147772 48188 147824
rect 18144 147704 18196 147756
rect 18696 147704 18748 147756
rect 58072 147704 58124 147756
rect 59360 147704 59412 147756
rect 18236 147636 18288 147688
rect 19248 147636 19300 147688
rect 19708 147636 19760 147688
rect 59544 147636 59596 147688
rect 19064 147568 19116 147620
rect 37004 147568 37056 147620
rect 48228 147568 48280 147620
rect 50160 147568 50212 147620
rect 63592 147568 63644 147620
rect 189724 147568 189776 147620
rect 406476 147568 406528 147620
rect 458364 147568 458416 147620
rect 459468 147568 459520 147620
rect 478052 147568 478104 147620
rect 16120 147500 16172 147552
rect 19340 147500 19392 147552
rect 20628 147500 20680 147552
rect 35900 147432 35952 147484
rect 19156 147364 19208 147416
rect 38108 147364 38160 147416
rect 18604 147296 18656 147348
rect 18972 147296 19024 147348
rect 19892 147296 19944 147348
rect 43076 147296 43128 147348
rect 61660 147500 61712 147552
rect 66168 147500 66220 147552
rect 180064 147500 180116 147552
rect 406660 147500 406712 147552
rect 455972 147500 456024 147552
rect 458088 147500 458140 147552
rect 476948 147500 477000 147552
rect 48136 147432 48188 147484
rect 51448 147432 51500 147484
rect 59544 147432 59596 147484
rect 78036 147432 78088 147484
rect 78496 147432 78548 147484
rect 188436 147432 188488 147484
rect 409144 147432 409196 147484
rect 453580 147432 453632 147484
rect 47676 147364 47728 147416
rect 66352 147364 66404 147416
rect 70400 147364 70452 147416
rect 75644 147364 75696 147416
rect 75828 147364 75880 147416
rect 79140 147364 79192 147416
rect 81072 147364 81124 147416
rect 188344 147364 188396 147416
rect 415124 147364 415176 147416
rect 448244 147364 448296 147416
rect 59360 147296 59412 147348
rect 76932 147296 76984 147348
rect 88248 147296 88300 147348
rect 186044 147296 186096 147348
rect 418344 147296 418396 147348
rect 450636 147296 450688 147348
rect 15660 147228 15712 147280
rect 19248 147228 19300 147280
rect 19800 147228 19852 147280
rect 44180 147228 44232 147280
rect 44732 147228 44784 147280
rect 46020 147228 46072 147280
rect 46572 147228 46624 147280
rect 65156 147228 65208 147280
rect 91008 147228 91060 147280
rect 185584 147228 185636 147280
rect 414664 147228 414716 147280
rect 440240 147228 440292 147280
rect 15936 147160 15988 147212
rect 16396 147160 16448 147212
rect 48688 147160 48740 147212
rect 67640 147160 67692 147212
rect 68284 147160 68336 147212
rect 162216 147160 162268 147212
rect 418712 147160 418764 147212
rect 419080 147160 419132 147212
rect 437020 147160 437072 147212
rect 18696 147092 18748 147144
rect 19156 147092 19208 147144
rect 19708 147092 19760 147144
rect 19892 147092 19944 147144
rect 21364 147092 21416 147144
rect 54024 147092 54076 147144
rect 71228 147092 71280 147144
rect 164056 147092 164108 147144
rect 419356 147092 419408 147144
rect 439596 147092 439648 147144
rect 16028 147024 16080 147076
rect 16488 147024 16540 147076
rect 52276 147024 52328 147076
rect 71044 147024 71096 147076
rect 95976 147024 96028 147076
rect 185768 147024 185820 147076
rect 419632 147024 419684 147076
rect 443092 147024 443144 147076
rect 461676 147024 461728 147076
rect 16304 146956 16356 147008
rect 53380 146956 53432 147008
rect 72148 146956 72200 147008
rect 103520 146956 103572 147008
rect 191104 146956 191156 147008
rect 418436 146956 418488 147008
rect 419264 146956 419316 147008
rect 444196 146956 444248 147008
rect 462780 146956 462832 147008
rect 18880 146888 18932 146940
rect 21364 146888 21416 146940
rect 18328 146820 18380 146872
rect 56048 146888 56100 146940
rect 73712 146888 73764 146940
rect 100944 146888 100996 146940
rect 182916 146888 182968 146940
rect 419724 146888 419776 146940
rect 419908 146888 419960 146940
rect 454592 146888 454644 146940
rect 473360 146888 473412 146940
rect 50160 146820 50212 146872
rect 68468 146820 68520 146872
rect 106096 146820 106148 146872
rect 156604 146820 156656 146872
rect 418620 146820 418672 146872
rect 419172 146820 419224 146872
rect 437940 146820 437992 146872
rect 445300 146820 445352 146872
rect 463884 146820 463936 146872
rect 51448 146752 51500 146804
rect 69756 146752 69808 146804
rect 108856 146752 108908 146804
rect 158168 146752 158220 146804
rect 418896 146752 418948 146804
rect 436100 146752 436152 146804
rect 447140 146752 447192 146804
rect 466276 146752 466328 146804
rect 18788 146480 18840 146532
rect 39580 146480 39632 146532
rect 18512 146412 18564 146464
rect 19248 146412 19300 146464
rect 45284 146684 45336 146736
rect 63868 146684 63920 146736
rect 111616 146684 111668 146736
rect 157984 146684 158036 146736
rect 430580 146684 430632 146736
rect 438216 146684 438268 146736
rect 448520 146684 448572 146736
rect 467564 146684 467616 146736
rect 44732 146616 44784 146668
rect 62764 146616 62816 146668
rect 449900 146616 449952 146668
rect 468668 146616 468720 146668
rect 54024 146548 54076 146600
rect 73252 146548 73304 146600
rect 452476 146548 452528 146600
rect 469772 146548 469824 146600
rect 452568 146480 452620 146532
rect 471060 146480 471112 146532
rect 446404 146412 446456 146464
rect 465172 146412 465224 146464
rect 15752 146344 15804 146396
rect 18604 146344 18656 146396
rect 46020 146344 46072 146396
rect 20628 146276 20680 146328
rect 47676 146276 47728 146328
rect 415768 146208 415820 146260
rect 416320 146208 416372 146260
rect 417148 146208 417200 146260
rect 417792 146208 417844 146260
rect 449900 146208 449952 146260
rect 419816 146140 419868 146192
rect 453396 146140 453448 146192
rect 472164 146344 472216 146396
rect 456800 146276 456852 146328
rect 474096 146276 474148 146328
rect 415676 146072 415728 146124
rect 416688 146072 416740 146124
rect 419448 146072 419500 146124
rect 452568 146072 452620 146124
rect 448520 146004 448572 146056
rect 419540 145936 419592 145988
rect 420000 145936 420052 145988
rect 451280 145936 451332 145988
rect 452476 145936 452528 145988
rect 416504 145868 416556 145920
rect 447140 145868 447192 145920
rect 417792 145800 417844 145852
rect 445300 145800 445352 145852
rect 418988 145732 419040 145784
rect 446404 145732 446456 145784
rect 531044 144848 531096 144900
rect 536840 144848 536892 144900
rect 577596 139340 577648 139392
rect 579620 139340 579672 139392
rect 536840 138660 536892 138712
rect 556896 138660 556948 138712
rect 3516 137912 3568 137964
rect 167828 137912 167880 137964
rect 151268 136552 151320 136604
rect 156696 136552 156748 136604
rect 551928 136552 551980 136604
rect 556804 136552 556856 136604
rect 418528 135192 418580 135244
rect 456800 135192 456852 135244
rect 187516 134648 187568 134700
rect 580448 134648 580500 134700
rect 187608 134580 187660 134632
rect 580908 134580 580960 134632
rect 187424 134512 187476 134564
rect 580356 134512 580408 134564
rect 417332 134376 417384 134428
rect 418528 134376 418580 134428
rect 3148 111732 3200 111784
rect 14740 111732 14792 111784
rect 556896 110372 556948 110424
rect 559564 110372 559616 110424
rect 577504 100648 577556 100700
rect 579712 100648 579764 100700
rect 559564 98948 559616 99000
rect 565084 98948 565136 99000
rect 3516 97928 3568 97980
rect 14648 97928 14700 97980
rect 565084 91740 565136 91792
rect 569960 91740 570012 91792
rect 161480 88952 161532 89004
rect 211160 88952 211212 89004
rect 269120 88952 269172 89004
rect 309784 88952 309836 89004
rect 267740 87592 267792 87644
rect 305644 87592 305696 87644
rect 233884 87320 233936 87372
rect 234620 87320 234672 87372
rect 190460 86232 190512 86284
rect 222200 86232 222252 86284
rect 302884 86232 302936 86284
rect 389180 86232 389232 86284
rect 3516 85484 3568 85536
rect 14556 85484 14608 85536
rect 569960 85484 570012 85536
rect 573364 85484 573416 85536
rect 573364 73108 573416 73160
rect 580172 73108 580224 73160
rect 3516 71680 3568 71732
rect 14464 71680 14516 71732
rect 393964 59304 394016 59356
rect 416780 59304 416832 59356
rect 418712 49920 418764 49972
rect 456984 49920 457036 49972
rect 16304 49852 16356 49904
rect 53472 49852 53524 49904
rect 417700 49852 417752 49904
rect 458088 49852 458140 49904
rect 17040 49784 17092 49836
rect 59544 49784 59596 49836
rect 408316 49784 408368 49836
rect 478512 49784 478564 49836
rect 15108 49716 15160 49768
rect 60648 49716 60700 49768
rect 408040 49716 408092 49768
rect 480904 49716 480956 49768
rect 95884 49648 95936 49700
rect 166632 49648 166684 49700
rect 407856 49648 407908 49700
rect 495900 49648 495952 49700
rect 91008 49580 91060 49632
rect 166448 49580 166500 49632
rect 413560 49580 413612 49632
rect 503536 49580 503588 49632
rect 88248 49512 88300 49564
rect 166540 49512 166592 49564
rect 410800 49512 410852 49564
rect 500960 49512 501012 49564
rect 86040 49444 86092 49496
rect 166816 49444 166868 49496
rect 406384 49444 406436 49496
rect 498476 49444 498528 49496
rect 83556 49376 83608 49428
rect 166356 49376 166408 49428
rect 410892 49376 410944 49428
rect 505928 49376 505980 49428
rect 80980 49308 81032 49360
rect 166724 49308 166776 49360
rect 413652 49308 413704 49360
rect 508504 49308 508556 49360
rect 58532 49240 58584 49292
rect 159640 49240 159692 49292
rect 413468 49240 413520 49292
rect 510988 49240 511040 49292
rect 56048 49172 56100 49224
rect 159732 49172 159784 49224
rect 416136 49172 416188 49224
rect 515864 49172 515916 49224
rect 53656 49104 53708 49156
rect 161204 49104 161256 49156
rect 413376 49104 413428 49156
rect 513380 49104 513432 49156
rect 50804 49036 50856 49088
rect 163872 49036 163924 49088
rect 411904 49036 411956 49088
rect 520924 49036 520976 49088
rect 48320 48968 48372 49020
rect 169300 48968 169352 49020
rect 416596 48968 416648 49020
rect 525892 48968 525944 49020
rect 98552 48900 98604 48952
rect 163688 48900 163740 48952
rect 410616 48900 410668 48952
rect 493416 48900 493468 48952
rect 103520 48832 103572 48884
rect 163964 48832 164016 48884
rect 407948 48832 408000 48884
rect 488264 48832 488316 48884
rect 106004 48764 106056 48816
rect 163780 48764 163832 48816
rect 418804 48764 418856 48816
rect 459928 48764 459980 48816
rect 19064 48220 19116 48272
rect 36820 48220 36872 48272
rect 59544 48220 59596 48272
rect 78036 48220 78088 48272
rect 125968 48220 126020 48272
rect 388076 48220 388128 48272
rect 416044 48220 416096 48272
rect 458364 48220 458416 48272
rect 459468 48220 459520 48272
rect 478052 48220 478104 48272
rect 19616 48152 19668 48204
rect 57060 48152 57112 48204
rect 61200 48152 61252 48204
rect 159364 48152 159416 48204
rect 405096 48152 405148 48204
rect 448244 48152 448296 48204
rect 458088 48152 458140 48204
rect 476948 48152 477000 48204
rect 18420 48084 18472 48136
rect 55864 48084 55916 48136
rect 56508 48084 56560 48136
rect 65984 48084 66036 48136
rect 161112 48084 161164 48136
rect 413284 48084 413336 48136
rect 453580 48084 453632 48136
rect 469128 48084 469180 48136
rect 475660 48084 475712 48136
rect 18880 48016 18932 48068
rect 16488 47948 16540 48000
rect 16396 47880 16448 47932
rect 48688 47880 48740 47932
rect 18144 47812 18196 47864
rect 51448 47812 51500 47864
rect 19984 47744 20036 47796
rect 49700 47744 49752 47796
rect 19340 47676 19392 47728
rect 47584 47676 47636 47728
rect 48228 47676 48280 47728
rect 63960 48016 64012 48068
rect 159548 48016 159600 48068
rect 410524 48016 410576 48068
rect 450636 48016 450688 48068
rect 53472 47948 53524 48000
rect 71780 47948 71832 48000
rect 73804 47948 73856 48000
rect 169116 47948 169168 48000
rect 417332 47948 417384 48000
rect 455880 47948 455932 48000
rect 474372 47948 474424 48000
rect 54576 47880 54628 47932
rect 73252 47880 73304 47932
rect 76104 47880 76156 47932
rect 169208 47880 169260 47932
rect 419724 47880 419776 47932
rect 454592 47880 454644 47932
rect 68376 47812 68428 47864
rect 159456 47812 159508 47864
rect 419264 47812 419316 47864
rect 444288 47812 444340 47864
rect 52368 47744 52420 47796
rect 71044 47744 71096 47796
rect 71136 47744 71188 47796
rect 162124 47744 162176 47796
rect 419632 47744 419684 47796
rect 67640 47676 67692 47728
rect 78496 47676 78548 47728
rect 169024 47676 169076 47728
rect 419356 47676 419408 47728
rect 439596 47676 439648 47728
rect 443092 47676 443144 47728
rect 461676 47676 461728 47728
rect 18604 47608 18656 47660
rect 46572 47608 46624 47660
rect 65064 47608 65116 47660
rect 93584 47608 93636 47660
rect 166264 47608 166316 47660
rect 419172 47608 419224 47660
rect 438124 47608 438176 47660
rect 444288 47608 444340 47660
rect 462780 47608 462832 47660
rect 18512 47540 18564 47592
rect 45376 47540 45428 47592
rect 19800 47472 19852 47524
rect 44180 47472 44232 47524
rect 48228 47540 48280 47592
rect 66260 47540 66312 47592
rect 100944 47540 100996 47592
rect 163596 47540 163648 47592
rect 418896 47540 418948 47592
rect 436100 47540 436152 47592
rect 473360 47540 473412 47592
rect 63868 47472 63920 47524
rect 111156 47472 111208 47524
rect 160744 47472 160796 47524
rect 419080 47472 419132 47524
rect 437020 47472 437072 47524
rect 19708 47404 19760 47456
rect 43168 47404 43220 47456
rect 61384 47404 61436 47456
rect 115848 47404 115900 47456
rect 160928 47404 160980 47456
rect 451280 47404 451332 47456
rect 469220 47404 469272 47456
rect 44180 47336 44232 47388
rect 62212 47336 62264 47388
rect 118608 47336 118660 47388
rect 160836 47336 160888 47388
rect 449532 47336 449584 47388
rect 467564 47336 467616 47388
rect 18236 47268 18288 47320
rect 57980 47268 58032 47320
rect 76380 47268 76432 47320
rect 450452 47268 450504 47320
rect 468668 47268 468720 47320
rect 50252 47200 50304 47252
rect 68560 47200 68612 47252
rect 447508 47200 447560 47252
rect 466276 47200 466328 47252
rect 56508 47132 56560 47184
rect 74356 47132 74408 47184
rect 451280 47132 451332 47184
rect 452292 47132 452344 47184
rect 471244 47132 471296 47184
rect 51448 47064 51500 47116
rect 69756 47064 69808 47116
rect 445300 47064 445352 47116
rect 463884 47064 463936 47116
rect 446404 46996 446456 47048
rect 465172 46996 465224 47048
rect 453948 46928 454000 46980
rect 472164 46928 472216 46980
rect 108856 46860 108908 46912
rect 163504 46860 163556 46912
rect 190276 46860 190328 46912
rect 580172 46860 580224 46912
rect 395344 46792 395396 46844
rect 470876 46792 470928 46844
rect 395528 46724 395580 46776
rect 468300 46724 468352 46776
rect 395436 46656 395488 46708
rect 465908 46656 465960 46708
rect 403624 46588 403676 46640
rect 463516 46588 463568 46640
rect 419816 46520 419868 46572
rect 453948 46520 454000 46572
rect 418988 46452 419040 46504
rect 446404 46452 446456 46504
rect 417792 46384 417844 46436
rect 445300 46384 445352 46436
rect 133880 46180 133932 46232
rect 199384 46180 199436 46232
rect 3424 45500 3476 45552
rect 167736 45500 167788 45552
rect 416320 45500 416372 45552
rect 450084 45500 450136 45552
rect 416688 45432 416740 45484
rect 449532 45432 449584 45484
rect 419448 45364 419500 45416
rect 451280 45364 451332 45416
rect 420000 45296 420052 45348
rect 451372 45296 451424 45348
rect 416504 45228 416556 45280
rect 447508 45228 447560 45280
rect 340880 44820 340932 44872
rect 494704 44820 494756 44872
rect 336740 43392 336792 43444
rect 483664 43392 483716 43444
rect 126980 42032 127032 42084
rect 197452 42032 197504 42084
rect 347780 42032 347832 42084
rect 512644 42032 512696 42084
rect 351920 40672 351972 40724
rect 523040 40672 523092 40724
rect 125600 39312 125652 39364
rect 194600 39312 194652 39364
rect 343640 39312 343692 39364
rect 502340 39312 502392 39364
rect 316040 37884 316092 37936
rect 431960 37884 432012 37936
rect 361580 36524 361632 36576
rect 547880 36524 547932 36576
rect 313924 35164 313976 35216
rect 420920 35164 420972 35216
rect 364340 33736 364392 33788
rect 555424 33736 555476 33788
rect 3148 33056 3200 33108
rect 167644 33056 167696 33108
rect 336004 32376 336056 32428
rect 473360 32376 473412 32428
rect 321560 31016 321612 31068
rect 445760 31016 445812 31068
rect 320180 29588 320232 29640
rect 441620 29588 441672 29640
rect 317420 28228 317472 28280
rect 434720 28228 434772 28280
rect 329104 26868 329156 26920
rect 456800 26868 456852 26920
rect 318800 25508 318852 25560
rect 438860 25508 438912 25560
rect 211160 24080 211212 24132
rect 230480 24080 230532 24132
rect 322940 24080 322992 24132
rect 448520 24080 448572 24132
rect 314660 22720 314712 22772
rect 427820 22720 427872 22772
rect 313280 21360 313332 21412
rect 423680 21360 423732 21412
rect 3424 20612 3476 20664
rect 170496 20612 170548 20664
rect 310520 17212 310572 17264
rect 416780 17212 416832 17264
rect 298744 15852 298796 15904
rect 364616 15852 364668 15904
rect 367100 15852 367152 15904
rect 563060 15852 563112 15904
rect 273260 14424 273312 14476
rect 322112 14424 322164 14476
rect 345020 14424 345072 14476
rect 506480 14424 506532 14476
rect 346400 13064 346452 13116
rect 508504 13064 508556 13116
rect 270500 11704 270552 11756
rect 314660 11704 314712 11756
rect 342260 11704 342312 11756
rect 498936 11704 498988 11756
rect 266360 10276 266412 10328
rect 303896 10276 303948 10328
rect 339500 10276 339552 10328
rect 492312 10276 492364 10328
rect 169576 8916 169628 8968
rect 213920 8916 213972 8968
rect 262220 8916 262272 8968
rect 291936 8916 291988 8968
rect 338120 8916 338172 8968
rect 488816 8916 488868 8968
rect 263600 7624 263652 7676
rect 294052 7624 294104 7676
rect 130568 7556 130620 7608
rect 198740 7556 198792 7608
rect 201500 7556 201552 7608
rect 226340 7556 226392 7608
rect 277400 7556 277452 7608
rect 332692 7556 332744 7608
rect 335360 7556 335412 7608
rect 481732 7556 481784 7608
rect 3424 6808 3476 6860
rect 170404 6808 170456 6860
rect 190368 6808 190420 6860
rect 580172 6808 580224 6860
rect 292580 6536 292632 6588
rect 371700 6536 371752 6588
rect 293960 6468 294012 6520
rect 375288 6468 375340 6520
rect 295340 6400 295392 6452
rect 378876 6400 378928 6452
rect 300860 6332 300912 6384
rect 393044 6332 393096 6384
rect 362960 6264 363012 6316
rect 552664 6264 552716 6316
rect 288440 6196 288492 6248
rect 361120 6196 361172 6248
rect 369860 6196 369912 6248
rect 570328 6196 570380 6248
rect 291200 6128 291252 6180
rect 368204 6128 368256 6180
rect 371240 6128 371292 6180
rect 573916 6128 573968 6180
rect 274640 5312 274692 5364
rect 325608 5312 325660 5364
rect 276020 5244 276072 5296
rect 329196 5244 329248 5296
rect 349160 5244 349212 5296
rect 517152 5244 517204 5296
rect 278780 5176 278832 5228
rect 336280 5176 336332 5228
rect 350540 5176 350592 5228
rect 520740 5176 520792 5228
rect 280160 5108 280212 5160
rect 339868 5108 339920 5160
rect 353300 5108 353352 5160
rect 527824 5108 527876 5160
rect 281540 5040 281592 5092
rect 343364 5040 343416 5092
rect 354680 5040 354732 5092
rect 531320 5040 531372 5092
rect 282920 4972 282972 5024
rect 346952 4972 347004 5024
rect 356060 4972 356112 5024
rect 534908 4972 534960 5024
rect 284300 4904 284352 4956
rect 350448 4904 350500 4956
rect 357440 4904 357492 4956
rect 538404 4904 538456 4956
rect 194416 4836 194468 4888
rect 223580 4836 223632 4888
rect 285680 4836 285732 4888
rect 354036 4836 354088 4888
rect 358820 4836 358872 4888
rect 541992 4836 542044 4888
rect 128176 4768 128228 4820
rect 195244 4768 195296 4820
rect 287060 4768 287112 4820
rect 357532 4768 357584 4820
rect 360200 4768 360252 4820
rect 545488 4768 545540 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 508504 4088 508556 4140
rect 510068 4088 510120 4140
rect 576124 4088 576176 4140
rect 577412 4088 577464 4140
rect 248420 3952 248472 4004
rect 258264 3952 258316 4004
rect 298100 3952 298152 4004
rect 385960 3952 386012 4004
rect 249800 3884 249852 3936
rect 261760 3884 261812 3936
rect 305000 3884 305052 3936
rect 403624 3884 403676 3936
rect 158904 3816 158956 3868
rect 209780 3816 209832 3868
rect 251180 3816 251232 3868
rect 265348 3816 265400 3868
rect 324320 3816 324372 3868
rect 453304 3816 453356 3868
rect 155408 3748 155460 3800
rect 208400 3748 208452 3800
rect 252560 3748 252612 3800
rect 268844 3748 268896 3800
rect 327080 3748 327132 3800
rect 460388 3748 460440 3800
rect 151820 3680 151872 3732
rect 207020 3680 207072 3732
rect 253940 3680 253992 3732
rect 272432 3680 272484 3732
rect 305644 3680 305696 3732
rect 307944 3680 307996 3732
rect 328460 3680 328512 3732
rect 463976 3680 464028 3732
rect 148324 3612 148376 3664
rect 205640 3612 205692 3664
rect 219256 3612 219308 3664
rect 224224 3612 224276 3664
rect 255320 3612 255372 3664
rect 276020 3612 276072 3664
rect 329840 3612 329892 3664
rect 467472 3612 467524 3664
rect 144736 3544 144788 3596
rect 204260 3544 204312 3596
rect 215668 3544 215720 3596
rect 222844 3544 222896 3596
rect 244280 3544 244332 3596
rect 247592 3544 247644 3596
rect 256700 3544 256752 3596
rect 279516 3544 279568 3596
rect 331220 3544 331272 3596
rect 471060 3544 471112 3596
rect 1676 3476 1728 3528
rect 15844 3476 15896 3528
rect 141240 3476 141292 3528
rect 202880 3476 202932 3528
rect 208584 3476 208636 3528
rect 220084 3476 220136 3528
rect 226340 3476 226392 3528
rect 228364 3476 228416 3528
rect 229836 3476 229888 3528
rect 237380 3476 237432 3528
rect 240508 3476 240560 3528
rect 241520 3476 241572 3528
rect 242900 3476 242952 3528
rect 244096 3476 244148 3528
rect 245660 3476 245712 3528
rect 251180 3476 251232 3528
rect 258080 3476 258132 3528
rect 283104 3476 283156 3528
rect 287704 3476 287756 3528
rect 290188 3476 290240 3528
rect 299480 3476 299532 3528
rect 300768 3476 300820 3528
rect 309784 3476 309836 3528
rect 311440 3476 311492 3528
rect 333980 3476 334032 3528
rect 478144 3476 478196 3528
rect 494704 3476 494756 3528
rect 495900 3476 495952 3528
rect 512644 3476 512696 3528
rect 513564 3476 513616 3528
rect 555424 3476 555476 3528
rect 556160 3476 556212 3528
rect 137652 3408 137704 3460
rect 201592 3408 201644 3460
rect 205088 3408 205140 3460
rect 218704 3408 218756 3460
rect 222752 3408 222804 3460
rect 233884 3408 233936 3460
rect 247040 3408 247092 3460
rect 254676 3408 254728 3460
rect 259460 3408 259512 3460
rect 286600 3408 286652 3460
rect 374000 3408 374052 3460
rect 581000 3408 581052 3460
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 233424 3204 233476 3256
rect 238760 3204 238812 3256
rect 578884 3204 578936 3256
rect 582196 3204 582248 3256
rect 237012 3000 237064 3052
rect 239404 3000 239456 3052
rect 291936 3000 291988 3052
rect 293684 3000 293736 3052
rect 294052 2864 294104 2916
rect 297272 2864 297324 2916
rect 483664 2864 483716 2916
rect 485228 2864 485280 2916
rect 558184 2864 558236 2916
rect 559748 2864 559800 2916
rect 562324 2864 562376 2916
rect 566832 2864 566884 2916
rect 423680 2728 423732 2780
rect 424968 2728 425020 2780
rect 448520 2728 448572 2780
rect 449808 2728 449860 2780
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 699718 8156 703520
rect 8116 699712 8168 699718
rect 8116 699654 8168 699660
rect 10324 699712 10376 699718
rect 10324 699654 10376 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 4804 632120 4856 632126
rect 2832 632088 2834 632097
rect 4804 632062 4856 632068
rect 2778 632023 2834 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3436 481030 3464 566879
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3528 482322 3556 514791
rect 3516 482316 3568 482322
rect 3516 482258 3568 482264
rect 3424 481024 3476 481030
rect 3424 480966 3476 480972
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 4816 464370 4844 632062
rect 7564 527196 7616 527202
rect 7564 527138 7616 527144
rect 7576 467158 7604 527138
rect 10336 468518 10364 699654
rect 23492 692102 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 23480 692096 23532 692102
rect 23480 692038 23532 692044
rect 40052 687954 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 690674 71820 702986
rect 89180 700330 89208 703520
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 71780 690668 71832 690674
rect 71780 690610 71832 690616
rect 40040 687948 40092 687954
rect 40040 687890 40092 687896
rect 104912 686526 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 689314 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700398 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 136640 689308 136692 689314
rect 136640 689250 136692 689256
rect 104900 686520 104952 686526
rect 104900 686462 104952 686468
rect 169772 685166 169800 702406
rect 202800 700398 202828 703520
rect 199384 700392 199436 700398
rect 199384 700334 199436 700340
rect 202788 700392 202840 700398
rect 202788 700334 202840 700340
rect 203524 700392 203576 700398
rect 203524 700334 203576 700340
rect 169760 685160 169812 685166
rect 169760 685102 169812 685108
rect 166448 684956 166500 684962
rect 166448 684898 166500 684904
rect 163964 684888 164016 684894
rect 163964 684830 164016 684836
rect 159272 684820 159324 684826
rect 159272 684762 159324 684768
rect 156880 684752 156932 684758
rect 156880 684694 156932 684700
rect 154304 684684 154356 684690
rect 154304 684626 154356 684632
rect 132960 684616 133012 684622
rect 132960 684558 133012 684564
rect 118608 684548 118660 684554
rect 118608 684490 118660 684496
rect 111064 683732 111116 683738
rect 111064 683674 111116 683680
rect 104256 683664 104308 683670
rect 104256 683606 104308 683612
rect 97080 683596 97132 683602
rect 97080 683538 97132 683544
rect 94688 683528 94740 683534
rect 94688 683470 94740 683476
rect 92296 683460 92348 683466
rect 92296 683402 92348 683408
rect 70768 683392 70820 683398
rect 70768 683334 70820 683340
rect 44180 683324 44232 683330
rect 44180 683266 44232 683272
rect 32496 683256 32548 683262
rect 32496 683198 32548 683204
rect 25320 681896 25372 681902
rect 25320 681838 25372 681844
rect 25332 679946 25360 681838
rect 27528 681828 27580 681834
rect 27528 681770 27580 681776
rect 27540 679946 27568 681770
rect 30102 680368 30158 680377
rect 30102 680303 30158 680312
rect 30116 679946 30144 680303
rect 32508 679946 32536 683198
rect 42064 682848 42116 682854
rect 42064 682790 42116 682796
rect 37188 681760 37240 681766
rect 37188 681702 37240 681708
rect 34886 680504 34942 680513
rect 34886 680439 34942 680448
rect 34900 679946 34928 680439
rect 37200 679946 37228 681702
rect 39672 680400 39724 680406
rect 39672 680342 39724 680348
rect 39684 679946 39712 680342
rect 42076 679946 42104 682790
rect 44088 682304 44140 682310
rect 44088 682246 44140 682252
rect 25024 679918 25360 679946
rect 27416 679918 27568 679946
rect 29808 679918 30144 679946
rect 32200 679918 32536 679946
rect 34592 679918 34928 679946
rect 36984 679918 37228 679946
rect 39376 679918 39712 679946
rect 41768 679918 42104 679946
rect 44100 679946 44128 682246
rect 44192 681766 44220 683266
rect 61200 682916 61252 682922
rect 61200 682858 61252 682864
rect 46846 682680 46902 682689
rect 46846 682615 46902 682624
rect 44180 681760 44232 681766
rect 44180 681702 44232 681708
rect 46860 679946 46888 682615
rect 53654 682408 53710 682417
rect 53654 682343 53710 682352
rect 51630 682272 51686 682281
rect 51630 682207 51686 682216
rect 49240 680468 49292 680474
rect 49240 680410 49292 680416
rect 49252 679946 49280 680410
rect 51644 679946 51672 682207
rect 44100 679918 44160 679946
rect 46552 679918 46888 679946
rect 48944 679918 49280 679946
rect 51336 679918 51672 679946
rect 53668 679810 53696 682343
rect 58808 682168 58860 682174
rect 58808 682110 58860 682116
rect 56416 680536 56468 680542
rect 56416 680478 56468 680484
rect 56428 679946 56456 680478
rect 58820 679946 58848 682110
rect 60740 681896 60792 681902
rect 60740 681838 60792 681844
rect 60752 681057 60780 681838
rect 60738 681048 60794 681057
rect 60738 680983 60794 680992
rect 61212 679946 61240 682858
rect 65984 682236 66036 682242
rect 65984 682178 66036 682184
rect 63408 682032 63460 682038
rect 63408 681974 63460 681980
rect 63420 679946 63448 681974
rect 65996 679946 66024 682178
rect 68376 680604 68428 680610
rect 68376 680546 68428 680552
rect 68388 679946 68416 680546
rect 70780 679946 70808 683334
rect 85120 682780 85172 682786
rect 85120 682722 85172 682728
rect 79968 682100 80020 682106
rect 79968 682042 80020 682048
rect 75550 682000 75606 682009
rect 75550 681935 75606 681944
rect 73068 681896 73120 681902
rect 73068 681838 73120 681844
rect 73080 679946 73108 681838
rect 75564 679946 75592 681935
rect 79048 681828 79100 681834
rect 79048 681770 79100 681776
rect 77944 680672 77996 680678
rect 77944 680614 77996 680620
rect 77956 679946 77984 680614
rect 56120 679918 56456 679946
rect 58512 679918 58848 679946
rect 60904 679918 61240 679946
rect 63296 679918 63448 679946
rect 65688 679918 66024 679946
rect 68080 679918 68416 679946
rect 70472 679918 70808 679946
rect 72864 679918 73108 679946
rect 75256 679918 75592 679946
rect 77648 679918 77984 679946
rect 53668 679782 53728 679810
rect 79060 679561 79088 681770
rect 79980 679946 80008 682042
rect 82728 680740 82780 680746
rect 82728 680682 82780 680688
rect 82740 679946 82768 680682
rect 85132 679946 85160 682722
rect 85488 681896 85540 681902
rect 85488 681838 85540 681844
rect 85500 681018 85528 681838
rect 87512 681760 87564 681766
rect 87512 681702 87564 681708
rect 85488 681012 85540 681018
rect 85488 680954 85540 680960
rect 87524 679946 87552 681702
rect 92308 679946 92336 683402
rect 94700 679946 94728 683470
rect 97092 679946 97120 683538
rect 99288 682712 99340 682718
rect 99288 682654 99340 682660
rect 98644 681760 98696 681766
rect 98644 681702 98696 681708
rect 79980 679918 80040 679946
rect 82432 679918 82768 679946
rect 84824 679918 85160 679946
rect 87216 679918 87552 679946
rect 92000 679918 92336 679946
rect 94392 679918 94728 679946
rect 96784 679918 97120 679946
rect 98656 679658 98684 681702
rect 99300 679946 99328 682654
rect 101864 682576 101916 682582
rect 101864 682518 101916 682524
rect 100760 682236 100812 682242
rect 100760 682178 100812 682184
rect 100772 681086 100800 682178
rect 100760 681080 100812 681086
rect 100760 681022 100812 681028
rect 101876 679946 101904 682518
rect 104268 679946 104296 683606
rect 111076 682718 111104 683674
rect 111064 682712 111116 682718
rect 111064 682654 111116 682660
rect 106648 682644 106700 682650
rect 106648 682586 106700 682592
rect 106660 679946 106688 682586
rect 108948 682508 109000 682514
rect 108948 682450 109000 682456
rect 107568 682168 107620 682174
rect 107568 682110 107620 682116
rect 107580 681154 107608 682110
rect 107568 681148 107620 681154
rect 107568 681090 107620 681096
rect 108960 679946 108988 682450
rect 111432 680808 111484 680814
rect 111432 680750 111484 680756
rect 111444 679946 111472 680750
rect 118620 679946 118648 684490
rect 130384 683868 130436 683874
rect 130384 683810 130436 683816
rect 124220 683800 124272 683806
rect 124220 683742 124272 683748
rect 124232 682582 124260 683742
rect 130396 682650 130424 683810
rect 130384 682644 130436 682650
rect 130384 682586 130436 682592
rect 124220 682576 124272 682582
rect 124220 682518 124272 682524
rect 130568 682372 130620 682378
rect 130568 682314 130620 682320
rect 128176 681896 128228 681902
rect 128176 681838 128228 681844
rect 125416 681828 125468 681834
rect 125416 681770 125468 681776
rect 123392 680876 123444 680882
rect 123392 680818 123444 680824
rect 123404 679946 123432 680818
rect 99176 679918 99328 679946
rect 101568 679918 101904 679946
rect 103960 679918 104296 679946
rect 106352 679918 106688 679946
rect 108744 679918 108988 679946
rect 111136 679918 111472 679946
rect 118312 679918 118648 679946
rect 123096 679918 123432 679946
rect 125428 679810 125456 681770
rect 128188 679946 128216 681838
rect 130580 679946 130608 682314
rect 132972 679946 133000 684558
rect 142160 684004 142212 684010
rect 142160 683946 142212 683952
rect 133880 683936 133932 683942
rect 133880 683878 133932 683884
rect 133892 682514 133920 683878
rect 142172 682854 142200 683946
rect 146944 682916 146996 682922
rect 146944 682858 146996 682864
rect 142160 682848 142212 682854
rect 142160 682790 142212 682796
rect 137284 682780 137336 682786
rect 137284 682722 137336 682728
rect 133880 682508 133932 682514
rect 133880 682450 133932 682456
rect 127880 679918 128216 679946
rect 130272 679918 130608 679946
rect 132664 679918 133000 679946
rect 125428 679782 125488 679810
rect 137296 679726 137324 682722
rect 144828 682508 144880 682514
rect 144828 682450 144880 682456
rect 142528 682440 142580 682446
rect 142528 682382 142580 682388
rect 140136 682168 140188 682174
rect 137742 682136 137798 682145
rect 140136 682110 140188 682116
rect 137742 682071 137798 682080
rect 137756 679946 137784 682071
rect 140148 679946 140176 682110
rect 142540 679946 142568 682382
rect 144276 682100 144328 682106
rect 144276 682042 144328 682048
rect 137448 679918 137784 679946
rect 139840 679918 140176 679946
rect 142232 679918 142568 679946
rect 137284 679720 137336 679726
rect 144288 679697 144316 682042
rect 144840 679946 144868 682450
rect 146956 681222 146984 682858
rect 149704 682576 149756 682582
rect 149704 682518 149756 682524
rect 147312 681964 147364 681970
rect 147312 681906 147364 681912
rect 146944 681216 146996 681222
rect 146944 681158 146996 681164
rect 147324 679946 147352 681906
rect 149716 679946 149744 682518
rect 154316 679946 154344 684626
rect 156892 679946 156920 684694
rect 159284 679946 159312 684762
rect 161388 684072 161440 684078
rect 161388 684014 161440 684020
rect 161400 680218 161428 684014
rect 144624 679918 144868 679946
rect 147016 679918 147352 679946
rect 149408 679918 149744 679946
rect 154192 679918 154344 679946
rect 156584 679918 156920 679946
rect 158976 679918 159312 679946
rect 161354 680190 161428 680218
rect 161354 679932 161382 680190
rect 163976 679946 164004 684830
rect 166460 679946 166488 684898
rect 171048 682644 171100 682650
rect 171048 682586 171100 682592
rect 168380 682304 168432 682310
rect 168380 682246 168432 682252
rect 168392 681358 168420 682246
rect 169760 682032 169812 682038
rect 169760 681974 169812 681980
rect 168838 681864 168894 681873
rect 168838 681799 168894 681808
rect 168380 681352 168432 681358
rect 168380 681294 168432 681300
rect 168852 679946 168880 681799
rect 163760 679918 164004 679946
rect 166152 679918 166488 679946
rect 168544 679918 168880 679946
rect 169772 679833 169800 681974
rect 169758 679824 169814 679833
rect 171060 679810 171088 682586
rect 198188 682576 198240 682582
rect 197174 682544 197230 682553
rect 198188 682518 198240 682524
rect 197174 682479 197230 682488
rect 185584 682304 185636 682310
rect 185584 682246 185636 682252
rect 183192 682236 183244 682242
rect 183192 682178 183244 682184
rect 173808 682168 173860 682174
rect 173808 682110 173860 682116
rect 178408 682168 178460 682174
rect 178408 682110 178460 682116
rect 173624 681760 173676 681766
rect 173624 681702 173676 681708
rect 173636 679946 173664 681702
rect 173820 681290 173848 682110
rect 176016 682032 176068 682038
rect 176016 681974 176068 681980
rect 173808 681284 173860 681290
rect 173808 681226 173860 681232
rect 176028 679946 176056 681974
rect 178420 679946 178448 682110
rect 180616 682100 180668 682106
rect 180616 682042 180668 682048
rect 180628 679946 180656 682042
rect 183204 679946 183232 682178
rect 185596 679946 185624 682246
rect 195150 682136 195206 682145
rect 195150 682071 195206 682080
rect 192758 682000 192814 682009
rect 192758 681935 192814 681944
rect 192772 679946 192800 681935
rect 195164 679946 195192 682071
rect 173328 679918 173664 679946
rect 175720 679918 176056 679946
rect 178112 679918 178448 679946
rect 180504 679918 180656 679946
rect 182896 679918 183232 679946
rect 185288 679918 185624 679946
rect 192464 679918 192800 679946
rect 194856 679918 195192 679946
rect 197188 679946 197216 682479
rect 198004 682440 198056 682446
rect 198004 682382 198056 682388
rect 197188 679918 197248 679946
rect 170936 679782 171088 679810
rect 169758 679759 169814 679768
rect 137284 679662 137336 679668
rect 144274 679688 144330 679697
rect 98644 679652 98696 679658
rect 144274 679623 144330 679632
rect 98644 679594 98696 679600
rect 79046 679552 79102 679561
rect 79046 679487 79102 679496
rect 89720 679448 89772 679454
rect 89608 679396 89720 679402
rect 113824 679448 113876 679454
rect 89608 679390 89772 679396
rect 113528 679396 113824 679402
rect 116032 679448 116084 679454
rect 113528 679390 113876 679396
rect 115920 679396 116032 679402
rect 121000 679448 121052 679454
rect 115920 679390 116084 679396
rect 120704 679396 121000 679402
rect 135168 679448 135220 679454
rect 120704 679390 121052 679396
rect 135056 679396 135168 679402
rect 151912 679448 151964 679454
rect 135056 679390 135220 679396
rect 151800 679396 151912 679402
rect 187792 679448 187844 679454
rect 151800 679390 151964 679396
rect 187680 679396 187792 679402
rect 187680 679390 187844 679396
rect 89608 679374 89760 679390
rect 113528 679374 113864 679390
rect 115920 679374 116072 679390
rect 120704 679374 121040 679390
rect 135056 679374 135208 679390
rect 151800 679374 151952 679390
rect 187680 679374 187832 679390
rect 190044 679280 190100 679289
rect 22112 679238 22632 679266
rect 20904 670744 20956 670750
rect 20904 670686 20956 670692
rect 20916 663794 20944 670686
rect 20916 663766 21404 663794
rect 11704 656940 11756 656946
rect 11704 656882 11756 656888
rect 11716 469878 11744 656882
rect 19984 618316 20036 618322
rect 19984 618258 20036 618264
rect 14464 605872 14516 605878
rect 14464 605814 14516 605820
rect 14476 471306 14504 605814
rect 18604 579692 18656 579698
rect 18604 579634 18656 579640
rect 15844 553444 15896 553450
rect 15844 553386 15896 553392
rect 15856 472666 15884 553386
rect 15844 472660 15896 472666
rect 15844 472602 15896 472608
rect 14464 471300 14516 471306
rect 14464 471242 14516 471248
rect 11704 469872 11756 469878
rect 11704 469814 11756 469820
rect 10324 468512 10376 468518
rect 10324 468454 10376 468460
rect 7564 467152 7616 467158
rect 7564 467094 7616 467100
rect 18616 465798 18644 579634
rect 19996 479602 20024 618258
rect 20076 501016 20128 501022
rect 20076 500958 20128 500964
rect 19984 479596 20036 479602
rect 19984 479538 20036 479544
rect 20088 474094 20116 500958
rect 21376 478174 21404 663766
rect 21364 478168 21416 478174
rect 21364 478110 21416 478116
rect 22112 476814 22140 679238
rect 190044 679215 190100 679224
rect 64952 500126 65288 500154
rect 65260 497486 65288 500126
rect 154592 500126 154928 500154
rect 65248 497480 65300 497486
rect 65248 497422 65300 497428
rect 151084 497480 151136 497486
rect 151084 497422 151136 497428
rect 22100 476808 22152 476814
rect 22100 476750 22152 476756
rect 20076 474088 20128 474094
rect 20076 474030 20128 474036
rect 18604 465792 18656 465798
rect 18604 465734 18656 465740
rect 14648 465248 14700 465254
rect 14648 465190 14700 465196
rect 4804 464364 4856 464370
rect 4804 464306 4856 464312
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 14556 462460 14608 462466
rect 14556 462402 14608 462408
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 14464 459808 14516 459814
rect 14464 459750 14516 459756
rect 4068 453008 4120 453014
rect 4068 452950 4120 452956
rect 3424 452940 3476 452946
rect 3424 452882 3476 452888
rect 3332 452872 3384 452878
rect 3332 452814 3384 452820
rect 3240 450628 3292 450634
rect 3240 450570 3292 450576
rect 3252 423609 3280 450570
rect 3238 423600 3294 423609
rect 3238 423535 3294 423544
rect 3344 410553 3372 452814
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3436 358465 3464 452882
rect 3606 452840 3662 452849
rect 3606 452775 3662 452784
rect 3792 452804 3844 452810
rect 3514 449576 3570 449585
rect 3514 449511 3516 449520
rect 3568 449511 3570 449520
rect 3516 449482 3568 449488
rect 3514 449440 3570 449449
rect 3514 449375 3570 449384
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3424 344344 3476 344350
rect 3424 344286 3476 344292
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 58585 3464 344286
rect 3528 254153 3556 449375
rect 3620 267209 3648 452775
rect 3792 452746 3844 452752
rect 3700 449744 3752 449750
rect 3700 449686 3752 449692
rect 3712 293185 3740 449686
rect 3804 306241 3832 452746
rect 3976 450016 4028 450022
rect 3976 449958 4028 449964
rect 3884 449676 3936 449682
rect 3884 449618 3936 449624
rect 3896 319297 3924 449618
rect 3988 371385 4016 449958
rect 4080 397497 4108 452950
rect 4066 397488 4122 397497
rect 4066 397423 4122 397432
rect 3974 371376 4030 371385
rect 3974 371311 4030 371320
rect 3882 319288 3938 319297
rect 3882 319223 3938 319232
rect 3790 306232 3846 306241
rect 3790 306167 3846 306176
rect 3698 293176 3754 293185
rect 3698 293111 3754 293120
rect 3606 267200 3662 267209
rect 3606 267135 3662 267144
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 7564 244928 7616 244934
rect 7564 244870 7616 244876
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 7576 4146 7604 244870
rect 14476 71738 14504 459750
rect 14568 85542 14596 462402
rect 14660 97986 14688 465190
rect 14924 459876 14976 459882
rect 14924 459818 14976 459824
rect 14832 454436 14884 454442
rect 14832 454378 14884 454384
rect 14738 449984 14794 449993
rect 14738 449919 14794 449928
rect 14752 111790 14780 449919
rect 14844 164218 14872 454378
rect 14936 189038 14964 459818
rect 15016 458244 15068 458250
rect 15016 458186 15068 458192
rect 15028 202842 15056 458186
rect 18972 455116 19024 455122
rect 18972 455058 19024 455064
rect 18880 454232 18932 454238
rect 18880 454174 18932 454180
rect 18788 454164 18840 454170
rect 18788 454106 18840 454112
rect 17408 453620 17460 453626
rect 17408 453562 17460 453568
rect 15106 452024 15162 452033
rect 15106 451959 15162 451968
rect 15120 215286 15148 451959
rect 17222 385928 17278 385937
rect 17222 385863 17278 385872
rect 16762 381032 16818 381041
rect 16762 380967 16818 380976
rect 16488 347268 16540 347274
rect 16488 347210 16540 347216
rect 16120 346792 16172 346798
rect 16120 346734 16172 346740
rect 16028 334620 16080 334626
rect 16028 334562 16080 334568
rect 15752 249076 15804 249082
rect 15752 249018 15804 249024
rect 15660 247648 15712 247654
rect 15660 247590 15712 247596
rect 15108 215280 15160 215286
rect 15108 215222 15160 215228
rect 15016 202836 15068 202842
rect 15016 202778 15068 202784
rect 14924 189032 14976 189038
rect 14924 188974 14976 188980
rect 14832 164212 14884 164218
rect 14832 164154 14884 164160
rect 15108 149116 15160 149122
rect 15108 149058 15160 149064
rect 14740 111784 14792 111790
rect 14740 111726 14792 111732
rect 14648 97980 14700 97986
rect 14648 97922 14700 97928
rect 14556 85536 14608 85542
rect 14556 85478 14608 85484
rect 14464 71732 14516 71738
rect 14464 71674 14516 71680
rect 15120 49774 15148 149058
rect 15672 147286 15700 247590
rect 15660 147280 15712 147286
rect 15660 147222 15712 147228
rect 15764 146402 15792 249018
rect 16040 247450 16068 334562
rect 16132 247858 16160 346734
rect 16212 346656 16264 346662
rect 16212 346598 16264 346604
rect 16120 247852 16172 247858
rect 16120 247794 16172 247800
rect 16028 247444 16080 247450
rect 16028 247386 16080 247392
rect 15936 247104 15988 247110
rect 15936 247046 15988 247052
rect 15844 233912 15896 233918
rect 15844 233854 15896 233860
rect 15752 146396 15804 146402
rect 15752 146338 15804 146344
rect 15108 49768 15160 49774
rect 15108 49710 15160 49716
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 584 480 612 4082
rect 15856 3534 15884 233854
rect 15948 147218 15976 247046
rect 16028 235748 16080 235754
rect 16028 235690 16080 235696
rect 15936 147212 15988 147218
rect 15936 147154 15988 147160
rect 16040 147082 16068 235690
rect 16132 147558 16160 247794
rect 16224 247790 16252 346598
rect 16304 346588 16356 346594
rect 16304 346530 16356 346536
rect 16316 248402 16344 346530
rect 16396 346520 16448 346526
rect 16396 346462 16448 346468
rect 16304 248396 16356 248402
rect 16304 248338 16356 248344
rect 16212 247784 16264 247790
rect 16212 247726 16264 247732
rect 16224 247110 16252 247726
rect 16212 247104 16264 247110
rect 16212 247046 16264 247052
rect 16304 235816 16356 235822
rect 16304 235758 16356 235764
rect 16120 147552 16172 147558
rect 16120 147494 16172 147500
rect 16028 147076 16080 147082
rect 16028 147018 16080 147024
rect 16316 147014 16344 235758
rect 16408 235754 16436 346462
rect 16500 235822 16528 347210
rect 16776 281081 16804 380967
rect 16946 359952 17002 359961
rect 16946 359887 17002 359896
rect 16854 283792 16910 283801
rect 16854 283727 16910 283736
rect 16762 281072 16818 281081
rect 16762 281007 16818 281016
rect 16488 235816 16540 235822
rect 16488 235758 16540 235764
rect 16396 235748 16448 235754
rect 16396 235690 16448 235696
rect 16762 186960 16818 186969
rect 16762 186895 16818 186904
rect 16396 147212 16448 147218
rect 16396 147154 16448 147160
rect 16304 147008 16356 147014
rect 16304 146950 16356 146956
rect 16316 49910 16344 146950
rect 16304 49904 16356 49910
rect 16304 49846 16356 49852
rect 16408 47938 16436 147154
rect 16488 147076 16540 147082
rect 16488 147018 16540 147024
rect 16500 48006 16528 147018
rect 16776 86873 16804 186895
rect 16868 183841 16896 283727
rect 16960 260817 16988 359887
rect 17038 358320 17094 358329
rect 17038 358255 17094 358264
rect 16946 260808 17002 260817
rect 16946 260743 17002 260752
rect 17052 259418 17080 358255
rect 17130 285832 17186 285841
rect 17130 285767 17186 285776
rect 17040 259412 17092 259418
rect 17040 259354 17092 259360
rect 17040 247444 17092 247450
rect 17040 247386 17092 247392
rect 16854 183832 16910 183841
rect 16854 183767 16910 183776
rect 16868 180794 16896 183767
rect 16868 180766 16988 180794
rect 16762 86864 16818 86873
rect 16762 86799 16818 86808
rect 16960 83745 16988 180766
rect 17052 147898 17080 247386
rect 17144 186969 17172 285767
rect 17236 285705 17264 385863
rect 17420 383654 17448 453562
rect 17776 453076 17828 453082
rect 17776 453018 17828 453024
rect 17590 386880 17646 386889
rect 17590 386815 17646 386824
rect 17500 384328 17552 384334
rect 17500 384270 17552 384276
rect 17328 383626 17448 383654
rect 17328 379953 17356 383626
rect 17314 379944 17370 379953
rect 17314 379879 17370 379888
rect 17222 285696 17278 285705
rect 17222 285631 17278 285640
rect 17328 279993 17356 379879
rect 17406 378176 17462 378185
rect 17406 378111 17462 378120
rect 17314 279984 17370 279993
rect 17314 279919 17370 279928
rect 17328 277394 17356 279919
rect 17420 278769 17448 378111
rect 17512 283801 17540 384270
rect 17604 286929 17632 386815
rect 17684 382288 17736 382294
rect 17684 382230 17736 382236
rect 17590 286920 17646 286929
rect 17590 286855 17646 286864
rect 17604 285841 17632 286855
rect 17590 285832 17646 285841
rect 17590 285767 17646 285776
rect 17498 283792 17554 283801
rect 17498 283727 17554 283736
rect 17590 282840 17646 282849
rect 17696 282826 17724 382230
rect 17788 378185 17816 453018
rect 17868 450560 17920 450566
rect 17868 450502 17920 450508
rect 17774 378176 17830 378185
rect 17774 378111 17830 378120
rect 17774 285696 17830 285705
rect 17774 285631 17830 285640
rect 17646 282798 17724 282826
rect 17590 282775 17646 282784
rect 17498 281072 17554 281081
rect 17498 281007 17554 281016
rect 17406 278760 17462 278769
rect 17406 278695 17462 278704
rect 17236 277366 17356 277394
rect 17130 186960 17186 186969
rect 17130 186895 17186 186904
rect 17130 186008 17186 186017
rect 17130 185943 17186 185952
rect 17040 147892 17092 147898
rect 17040 147834 17092 147840
rect 16946 83736 17002 83745
rect 16946 83671 17002 83680
rect 17052 49842 17080 147834
rect 17144 85921 17172 185943
rect 17236 179489 17264 277366
rect 17406 260808 17462 260817
rect 17406 260743 17462 260752
rect 17420 260001 17448 260743
rect 17406 259992 17462 260001
rect 17406 259927 17462 259936
rect 17316 259412 17368 259418
rect 17316 259354 17368 259360
rect 17328 258369 17356 259354
rect 17314 258360 17370 258369
rect 17314 258295 17370 258304
rect 17328 235958 17356 258295
rect 17316 235952 17368 235958
rect 17316 235894 17368 235900
rect 17222 179480 17278 179489
rect 17222 179415 17278 179424
rect 17328 158409 17356 235894
rect 17420 160041 17448 259927
rect 17512 181121 17540 281007
rect 17604 182889 17632 282775
rect 17682 278760 17738 278769
rect 17682 278695 17738 278704
rect 17696 278225 17724 278695
rect 17682 278216 17738 278225
rect 17682 278151 17738 278160
rect 17590 182880 17646 182889
rect 17590 182815 17646 182824
rect 17498 181112 17554 181121
rect 17498 181047 17554 181056
rect 17406 160032 17462 160041
rect 17406 159967 17462 159976
rect 17314 158400 17370 158409
rect 17314 158335 17370 158344
rect 17130 85912 17186 85921
rect 17130 85847 17186 85856
rect 17328 58313 17356 158335
rect 17420 59945 17448 159967
rect 17512 81025 17540 181047
rect 17604 82929 17632 182815
rect 17696 180794 17724 278151
rect 17788 186017 17816 285631
rect 17880 258233 17908 450502
rect 18800 385937 18828 454106
rect 18786 385928 18842 385937
rect 18786 385863 18842 385872
rect 18892 384334 18920 454174
rect 18880 384328 18932 384334
rect 18880 384270 18932 384276
rect 18892 383761 18920 384270
rect 18878 383752 18934 383761
rect 18878 383687 18934 383696
rect 18984 382809 19012 455058
rect 19064 455048 19116 455054
rect 19064 454990 19116 454996
rect 18970 382800 19026 382809
rect 18970 382735 19026 382744
rect 18984 382294 19012 382735
rect 18972 382288 19024 382294
rect 18972 382230 19024 382236
rect 19076 381041 19104 454990
rect 19340 454096 19392 454102
rect 19340 454038 19392 454044
rect 19248 449948 19300 449954
rect 19248 449890 19300 449896
rect 19156 434036 19208 434042
rect 19156 433978 19208 433984
rect 19062 381032 19118 381041
rect 19062 380967 19118 380976
rect 19168 359961 19196 433978
rect 19154 359952 19210 359961
rect 19154 359887 19210 359896
rect 19260 358057 19288 449890
rect 19352 386889 19380 454038
rect 134338 449712 134394 449721
rect 134338 449647 134394 449656
rect 134352 444786 134380 449647
rect 131764 444780 131816 444786
rect 131764 444722 131816 444728
rect 134340 444780 134392 444786
rect 134340 444722 134392 444728
rect 131776 434042 131804 444722
rect 151096 435402 151124 497422
rect 151084 435396 151136 435402
rect 151084 435338 151136 435344
rect 151096 435305 151124 435338
rect 151082 435296 151138 435305
rect 151082 435231 151138 435240
rect 154592 434042 154620 500126
rect 197636 466608 197688 466614
rect 197636 466550 197688 466556
rect 196072 466540 196124 466546
rect 196072 466482 196124 466488
rect 160744 465520 160796 465526
rect 160744 465462 160796 465468
rect 159732 463208 159784 463214
rect 159732 463150 159784 463156
rect 159640 463140 159692 463146
rect 159640 463082 159692 463088
rect 159364 463072 159416 463078
rect 159364 463014 159416 463020
rect 156696 459672 156748 459678
rect 156696 459614 156748 459620
rect 156602 450120 156658 450129
rect 156602 450055 156658 450064
rect 131764 434036 131816 434042
rect 131764 433978 131816 433984
rect 154580 434036 154632 434042
rect 154580 433978 154632 433984
rect 19338 386880 19394 386889
rect 19338 386815 19394 386824
rect 19246 358048 19302 358057
rect 19246 357983 19302 357992
rect 91006 349888 91062 349897
rect 91006 349823 91062 349832
rect 93490 349888 93546 349897
rect 93490 349823 93546 349832
rect 98550 349888 98606 349897
rect 98550 349823 98606 349832
rect 103518 349888 103574 349897
rect 103518 349823 103574 349832
rect 38474 349616 38530 349625
rect 38474 349551 38530 349560
rect 50802 349616 50858 349625
rect 50802 349551 50858 349560
rect 56046 349616 56102 349625
rect 56046 349551 56102 349560
rect 58530 349616 58586 349625
rect 58530 349551 58586 349560
rect 61106 349616 61162 349625
rect 61106 349551 61162 349560
rect 62854 349616 62910 349625
rect 62854 349551 62910 349560
rect 68742 349616 68798 349625
rect 68742 349551 68798 349560
rect 72238 349616 72294 349625
rect 72238 349551 72294 349560
rect 38488 348634 38516 349551
rect 50816 348770 50844 349551
rect 53654 349072 53710 349081
rect 53654 349007 53710 349016
rect 50804 348764 50856 348770
rect 50804 348706 50856 348712
rect 39580 348696 39632 348702
rect 39580 348638 39632 348644
rect 38476 348628 38528 348634
rect 38476 348570 38528 348576
rect 38488 347886 38516 348570
rect 19156 347880 19208 347886
rect 19156 347822 19208 347828
rect 38476 347880 38528 347886
rect 38476 347822 38528 347828
rect 18696 347812 18748 347818
rect 18696 347754 18748 347760
rect 18604 346860 18656 346866
rect 18604 346802 18656 346808
rect 18236 346724 18288 346730
rect 18236 346666 18288 346672
rect 17866 258224 17922 258233
rect 17866 258159 17922 258168
rect 18248 235618 18276 346666
rect 18328 334892 18380 334898
rect 18328 334834 18380 334840
rect 18340 235890 18368 334834
rect 18512 334756 18564 334762
rect 18512 334698 18564 334704
rect 18524 247722 18552 334698
rect 18616 249082 18644 346802
rect 18708 249801 18736 347754
rect 18972 346928 19024 346934
rect 18972 346870 19024 346876
rect 18880 334960 18932 334966
rect 18880 334902 18932 334908
rect 18788 334824 18840 334830
rect 18788 334766 18840 334772
rect 18694 249792 18750 249801
rect 18694 249727 18750 249736
rect 18604 249076 18656 249082
rect 18604 249018 18656 249024
rect 18604 248260 18656 248266
rect 18604 248202 18656 248208
rect 18512 247716 18564 247722
rect 18512 247658 18564 247664
rect 18524 247178 18552 247658
rect 18512 247172 18564 247178
rect 18512 247114 18564 247120
rect 18328 235884 18380 235890
rect 18328 235826 18380 235832
rect 18236 235612 18288 235618
rect 18236 235554 18288 235560
rect 18248 235142 18276 235554
rect 18236 235136 18288 235142
rect 18236 235078 18288 235084
rect 17774 186008 17830 186017
rect 17774 185943 17830 185952
rect 17696 180766 17816 180794
rect 17788 178265 17816 180766
rect 17866 180024 17922 180033
rect 17866 179959 17922 179968
rect 17880 179489 17908 179959
rect 17866 179480 17922 179489
rect 17866 179415 17922 179424
rect 17774 178256 17830 178265
rect 17774 178191 17830 178200
rect 17590 82920 17646 82929
rect 17590 82855 17646 82864
rect 17498 81016 17554 81025
rect 17498 80951 17554 80960
rect 17788 78169 17816 178191
rect 17880 79937 17908 179415
rect 18144 147756 18196 147762
rect 18144 147698 18196 147704
rect 17866 79928 17922 79937
rect 17866 79863 17922 79872
rect 17774 78160 17830 78169
rect 17774 78095 17830 78104
rect 17406 59936 17462 59945
rect 17406 59871 17462 59880
rect 17314 58304 17370 58313
rect 17314 58239 17370 58248
rect 17040 49836 17092 49842
rect 17040 49778 17092 49784
rect 16488 48000 16540 48006
rect 16488 47942 16540 47948
rect 16396 47932 16448 47938
rect 16396 47874 16448 47880
rect 18156 47870 18184 147698
rect 18236 147688 18288 147694
rect 18236 147630 18288 147636
rect 18144 47864 18196 47870
rect 18144 47806 18196 47812
rect 18248 47326 18276 147630
rect 18340 146878 18368 235826
rect 18616 147354 18644 248202
rect 18696 235136 18748 235142
rect 18696 235078 18748 235084
rect 18708 147762 18736 235078
rect 18800 235006 18828 334766
rect 18892 235686 18920 334902
rect 18984 247654 19012 346870
rect 19168 248130 19196 347822
rect 39592 347818 39620 348638
rect 53668 348430 53696 349007
rect 56060 348906 56088 349551
rect 58544 348974 58572 349551
rect 61120 349042 61148 349551
rect 62868 349178 62896 349551
rect 68756 349246 68784 349551
rect 72252 349314 72280 349551
rect 91020 349450 91048 349823
rect 93504 349518 93532 349823
rect 98564 349586 98592 349823
rect 103532 349654 103560 349823
rect 103520 349648 103572 349654
rect 103520 349590 103572 349596
rect 98552 349580 98604 349586
rect 98552 349522 98604 349528
rect 93492 349512 93544 349518
rect 93492 349454 93544 349460
rect 91008 349444 91060 349450
rect 91008 349386 91060 349392
rect 78036 349376 78088 349382
rect 78036 349318 78088 349324
rect 71780 349308 71832 349314
rect 71780 349250 71832 349256
rect 72240 349308 72292 349314
rect 72240 349250 72292 349256
rect 67640 349240 67692 349246
rect 67640 349182 67692 349188
rect 68744 349240 68796 349246
rect 68744 349182 68796 349188
rect 62856 349172 62908 349178
rect 62856 349114 62908 349120
rect 62028 349104 62080 349110
rect 62026 349072 62028 349081
rect 62080 349072 62082 349081
rect 61108 349036 61160 349042
rect 62026 349007 62082 349016
rect 61108 348978 61160 348984
rect 58532 348968 58584 348974
rect 58532 348910 58584 348916
rect 56048 348900 56100 348906
rect 56048 348842 56100 348848
rect 53656 348424 53708 348430
rect 53656 348366 53708 348372
rect 39580 347812 39632 347818
rect 39580 347754 39632 347760
rect 39592 347721 39620 347754
rect 62040 347750 62068 349007
rect 42800 347744 42852 347750
rect 36174 347712 36230 347721
rect 36174 347647 36230 347656
rect 39578 347712 39634 347721
rect 39578 347647 39634 347656
rect 42798 347712 42800 347721
rect 62028 347744 62080 347750
rect 42852 347712 42854 347721
rect 42798 347647 42854 347656
rect 44178 347712 44234 347721
rect 44178 347647 44234 347656
rect 45374 347712 45430 347721
rect 46570 347712 46626 347721
rect 45374 347647 45430 347656
rect 45928 347676 45980 347682
rect 19616 347132 19668 347138
rect 19616 347074 19668 347080
rect 19524 334688 19576 334694
rect 19524 334630 19576 334636
rect 19340 249756 19392 249762
rect 19340 249698 19392 249704
rect 19352 248414 19380 249698
rect 19432 249620 19484 249626
rect 19432 249562 19484 249568
rect 19260 248386 19380 248414
rect 19260 248334 19288 248386
rect 19248 248328 19300 248334
rect 19248 248270 19300 248276
rect 19156 248124 19208 248130
rect 19156 248066 19208 248072
rect 18972 247648 19024 247654
rect 18972 247590 19024 247596
rect 19064 247104 19116 247110
rect 19064 247046 19116 247052
rect 18880 235680 18932 235686
rect 18880 235622 18932 235628
rect 18788 235000 18840 235006
rect 18788 234942 18840 234948
rect 18696 147756 18748 147762
rect 18696 147698 18748 147704
rect 18604 147348 18656 147354
rect 18604 147290 18656 147296
rect 18696 147144 18748 147150
rect 18696 147086 18748 147092
rect 18328 146872 18380 146878
rect 18328 146814 18380 146820
rect 18340 142154 18368 146814
rect 18512 146464 18564 146470
rect 18512 146406 18564 146412
rect 18340 142126 18460 142154
rect 18432 48142 18460 142126
rect 18420 48136 18472 48142
rect 18420 48078 18472 48084
rect 18524 47598 18552 146406
rect 18604 146396 18656 146402
rect 18604 146338 18656 146344
rect 18616 47666 18644 146338
rect 18708 47841 18736 147086
rect 18892 146946 18920 235622
rect 19076 147626 19104 247046
rect 19064 147620 19116 147626
rect 19064 147562 19116 147568
rect 18972 147348 19024 147354
rect 18972 147290 19024 147296
rect 18880 146940 18932 146946
rect 18880 146882 18932 146888
rect 18786 146840 18842 146849
rect 18786 146775 18842 146784
rect 18800 146538 18828 146775
rect 18788 146532 18840 146538
rect 18788 146474 18840 146480
rect 18800 47977 18828 146474
rect 18892 48074 18920 146882
rect 18880 48068 18932 48074
rect 18880 48010 18932 48016
rect 18786 47968 18842 47977
rect 18786 47903 18842 47912
rect 18694 47832 18750 47841
rect 18694 47767 18750 47776
rect 18604 47660 18656 47666
rect 18604 47602 18656 47608
rect 18512 47592 18564 47598
rect 18984 47569 19012 147290
rect 19076 48278 19104 147562
rect 19168 147422 19196 248066
rect 19260 247110 19288 248270
rect 19444 248266 19472 249562
rect 19536 248414 19564 334630
rect 19628 249762 19656 347074
rect 19892 347064 19944 347070
rect 19892 347006 19944 347012
rect 19800 346996 19852 347002
rect 19800 346938 19852 346944
rect 19708 346452 19760 346458
rect 19708 346394 19760 346400
rect 19616 249756 19668 249762
rect 19616 249698 19668 249704
rect 19720 249626 19748 346394
rect 19708 249620 19760 249626
rect 19708 249562 19760 249568
rect 19708 248464 19760 248470
rect 19536 248386 19656 248414
rect 19708 248406 19760 248412
rect 19432 248260 19484 248266
rect 19432 248202 19484 248208
rect 19628 248033 19656 248386
rect 19614 248024 19670 248033
rect 19614 247959 19670 247968
rect 19340 247172 19392 247178
rect 19340 247114 19392 247120
rect 19248 247104 19300 247110
rect 19248 247046 19300 247052
rect 19352 246922 19380 247114
rect 19432 247104 19484 247110
rect 19432 247046 19484 247052
rect 19260 246894 19380 246922
rect 19260 147694 19288 246894
rect 19248 147688 19300 147694
rect 19248 147630 19300 147636
rect 19340 147552 19392 147558
rect 19340 147494 19392 147500
rect 19156 147416 19208 147422
rect 19156 147358 19208 147364
rect 19168 147150 19196 147358
rect 19248 147280 19300 147286
rect 19248 147222 19300 147228
rect 19156 147144 19208 147150
rect 19156 147086 19208 147092
rect 19260 146470 19288 147222
rect 19248 146464 19300 146470
rect 19248 146406 19300 146412
rect 19064 48272 19116 48278
rect 19064 48214 19116 48220
rect 19352 47734 19380 147494
rect 19444 147393 19472 247046
rect 19524 235272 19576 235278
rect 19524 235214 19576 235220
rect 19536 235006 19564 235214
rect 19524 235000 19576 235006
rect 19524 234942 19576 234948
rect 19430 147384 19486 147393
rect 19430 147319 19486 147328
rect 19444 142154 19472 147319
rect 19536 147257 19564 234942
rect 19628 149122 19656 247959
rect 19616 149116 19668 149122
rect 19616 149058 19668 149064
rect 19628 148714 19656 149058
rect 19616 148708 19668 148714
rect 19616 148650 19668 148656
rect 19720 148442 19748 248406
rect 19812 247926 19840 346938
rect 19904 247994 19932 347006
rect 36188 346390 36216 347647
rect 37186 347304 37242 347313
rect 37186 347239 37242 347248
rect 37200 347138 37228 347239
rect 37188 347132 37240 347138
rect 37188 347074 37240 347080
rect 42812 347070 42840 347647
rect 44192 347614 44220 347647
rect 44180 347608 44232 347614
rect 44180 347550 44232 347556
rect 42800 347064 42852 347070
rect 42800 347006 42852 347012
rect 44192 347002 44220 347550
rect 45388 347206 45416 347647
rect 46570 347647 46572 347656
rect 45928 347618 45980 347624
rect 46624 347647 46626 347656
rect 47582 347712 47638 347721
rect 47582 347647 47638 347656
rect 48594 347712 48650 347721
rect 48594 347647 48650 347656
rect 50066 347712 50122 347721
rect 50066 347647 50122 347656
rect 51262 347712 51318 347721
rect 51262 347647 51318 347656
rect 52366 347712 52422 347721
rect 52366 347647 52422 347656
rect 53470 347712 53526 347721
rect 62028 347686 62080 347692
rect 53470 347647 53526 347656
rect 46572 347618 46624 347624
rect 45376 347200 45428 347206
rect 45376 347142 45428 347148
rect 44180 346996 44232 347002
rect 44180 346938 44232 346944
rect 41786 346896 41842 346905
rect 45940 346866 45968 347618
rect 41786 346831 41842 346840
rect 45928 346860 45980 346866
rect 41326 346488 41382 346497
rect 41326 346423 41382 346432
rect 36176 346384 36228 346390
rect 36176 346326 36228 346332
rect 41340 345098 41368 346423
rect 41800 345273 41828 346831
rect 45928 346802 45980 346808
rect 47596 346798 47624 347647
rect 47584 346792 47636 346798
rect 47584 346734 47636 346740
rect 48608 346662 48636 347647
rect 50080 347410 50108 347647
rect 51080 347540 51132 347546
rect 51080 347482 51132 347488
rect 50068 347404 50120 347410
rect 50068 347346 50120 347352
rect 49608 347132 49660 347138
rect 49608 347074 49660 347080
rect 49620 346662 49648 347074
rect 48596 346656 48648 346662
rect 48596 346598 48648 346604
rect 49608 346656 49660 346662
rect 49608 346598 49660 346604
rect 50080 346594 50108 347346
rect 50068 346588 50120 346594
rect 50068 346530 50120 346536
rect 51092 346526 51120 347482
rect 51276 346594 51304 347647
rect 52380 347546 52408 347647
rect 52368 347540 52420 347546
rect 52368 347482 52420 347488
rect 53484 347478 53512 347647
rect 62868 347614 62896 349114
rect 65156 348492 65208 348498
rect 65156 348434 65208 348440
rect 64788 347744 64840 347750
rect 63682 347712 63738 347721
rect 63682 347647 63738 347656
rect 64786 347712 64788 347721
rect 65168 347721 65196 348434
rect 64840 347712 64842 347721
rect 64786 347647 64842 347656
rect 65154 347712 65210 347721
rect 65154 347647 65156 347656
rect 62856 347608 62908 347614
rect 62856 347550 62908 347556
rect 53472 347472 53524 347478
rect 53472 347414 53524 347420
rect 56598 347440 56654 347449
rect 56598 347375 56654 347384
rect 59358 347440 59414 347449
rect 59358 347375 59414 347384
rect 60830 347440 60886 347449
rect 60830 347375 60886 347384
rect 56612 347274 56640 347375
rect 56600 347268 56652 347274
rect 56600 347210 56652 347216
rect 55126 346760 55182 346769
rect 55182 346730 55260 346746
rect 55182 346724 55272 346730
rect 55182 346718 55220 346724
rect 55126 346695 55182 346704
rect 55220 346666 55272 346672
rect 51264 346588 51316 346594
rect 51264 346530 51316 346536
rect 51080 346520 51132 346526
rect 51080 346462 51132 346468
rect 41786 345264 41842 345273
rect 41786 345199 41842 345208
rect 42706 345264 42762 345273
rect 42706 345199 42762 345208
rect 19984 345092 20036 345098
rect 19984 345034 20036 345040
rect 41328 345092 41380 345098
rect 41328 345034 41380 345040
rect 19996 248062 20024 345034
rect 42720 345030 42748 345199
rect 42708 345024 42760 345030
rect 42708 344966 42760 344972
rect 55232 334966 55260 346666
rect 55220 334960 55272 334966
rect 55220 334902 55272 334908
rect 56612 334898 56640 347210
rect 57978 347168 58034 347177
rect 57978 347103 58034 347112
rect 57992 346497 58020 347103
rect 59372 346662 59400 347375
rect 60738 347168 60794 347177
rect 60738 347103 60794 347112
rect 59360 346656 59412 346662
rect 59360 346598 59412 346604
rect 57978 346488 58034 346497
rect 57978 346423 58034 346432
rect 56600 334892 56652 334898
rect 56600 334834 56652 334840
rect 57992 334830 58020 346423
rect 57980 334824 58032 334830
rect 57980 334766 58032 334772
rect 59372 334762 59400 346598
rect 59360 334756 59412 334762
rect 59360 334698 59412 334704
rect 60752 334694 60780 347103
rect 60844 347002 60872 347375
rect 61934 347168 61990 347177
rect 61934 347103 61990 347112
rect 60832 346996 60884 347002
rect 60832 346938 60884 346944
rect 60740 334688 60792 334694
rect 60740 334630 60792 334636
rect 60844 334626 60872 346938
rect 61948 346526 61976 347103
rect 61936 346520 61988 346526
rect 61936 346462 61988 346468
rect 63696 346322 63724 347647
rect 64800 347206 64828 347647
rect 65208 347647 65210 347656
rect 65982 347712 66038 347721
rect 65982 347647 66038 347656
rect 66258 347712 66314 347721
rect 66258 347647 66260 347656
rect 65156 347618 65208 347624
rect 64788 347200 64840 347206
rect 64788 347142 64840 347148
rect 63684 346316 63736 346322
rect 63684 346258 63736 346264
rect 65996 346254 66024 347647
rect 66312 347647 66314 347656
rect 66260 347618 66312 347624
rect 66272 347070 66300 347618
rect 67652 347410 67680 349182
rect 68374 349072 68430 349081
rect 68374 349007 68430 349016
rect 68388 348294 68416 349007
rect 71136 348560 71188 348566
rect 71136 348502 71188 348508
rect 68376 348288 68428 348294
rect 68376 348230 68428 348236
rect 71148 347721 71176 348502
rect 67730 347712 67786 347721
rect 67730 347647 67786 347656
rect 71134 347712 71190 347721
rect 71134 347647 71190 347656
rect 67744 347614 67772 347647
rect 67732 347608 67784 347614
rect 67732 347550 67784 347556
rect 67640 347404 67692 347410
rect 67640 347346 67692 347352
rect 67744 347138 67772 347550
rect 71148 347546 71176 347647
rect 71136 347540 71188 347546
rect 71136 347482 71188 347488
rect 71792 347478 71820 349250
rect 74354 348528 74410 348537
rect 74354 348463 74410 348472
rect 74368 348226 74396 348463
rect 73160 348220 73212 348226
rect 73160 348162 73212 348168
rect 74356 348220 74408 348226
rect 74356 348162 74408 348168
rect 71780 347472 71832 347478
rect 71780 347414 71832 347420
rect 73172 347274 73200 348162
rect 78048 347721 78076 349318
rect 78494 349072 78550 349081
rect 78494 349007 78550 349016
rect 86038 349072 86094 349081
rect 86038 349007 86094 349016
rect 78508 348838 78536 349007
rect 78496 348832 78548 348838
rect 78496 348774 78548 348780
rect 86052 348362 86080 349007
rect 86040 348356 86092 348362
rect 86040 348298 86092 348304
rect 73250 347712 73306 347721
rect 73250 347647 73306 347656
rect 73710 347712 73766 347721
rect 73710 347647 73766 347656
rect 75458 347712 75514 347721
rect 75458 347647 75514 347656
rect 76102 347712 76158 347721
rect 76102 347647 76158 347656
rect 76746 347712 76802 347721
rect 76746 347647 76802 347656
rect 78034 347712 78090 347721
rect 78034 347647 78090 347656
rect 79138 347712 79194 347721
rect 79138 347647 79194 347656
rect 81070 347712 81126 347721
rect 81070 347647 81126 347656
rect 83646 347712 83702 347721
rect 83646 347647 83702 347656
rect 96066 347712 96122 347721
rect 96066 347647 96122 347656
rect 100942 347712 100998 347721
rect 100942 347647 100998 347656
rect 106094 347712 106150 347721
rect 106094 347647 106150 347656
rect 108670 347712 108726 347721
rect 108670 347647 108726 347656
rect 111062 347712 111118 347721
rect 111062 347647 111118 347656
rect 113454 347712 113510 347721
rect 113454 347647 113510 347656
rect 115846 347712 115902 347721
rect 115846 347647 115902 347656
rect 118606 347712 118662 347721
rect 118606 347647 118662 347656
rect 120998 347712 121054 347721
rect 120998 347647 121054 347656
rect 123390 347712 123446 347721
rect 123390 347647 123446 347656
rect 125966 347712 126022 347721
rect 125966 347647 126022 347656
rect 73264 347546 73292 347647
rect 73252 347540 73304 347546
rect 73252 347482 73304 347488
rect 73160 347268 73212 347274
rect 73160 347210 73212 347216
rect 69294 347168 69350 347177
rect 67732 347132 67784 347138
rect 69294 347103 69350 347112
rect 67732 347074 67784 347080
rect 66260 347064 66312 347070
rect 66260 347006 66312 347012
rect 69308 346594 69336 347103
rect 73264 346730 73292 347482
rect 73724 347342 73752 347647
rect 73712 347336 73764 347342
rect 73712 347278 73764 347284
rect 75472 347070 75500 347647
rect 76116 347410 76144 347647
rect 76760 347478 76788 347647
rect 76748 347472 76800 347478
rect 76748 347414 76800 347420
rect 76104 347404 76156 347410
rect 76104 347346 76156 347352
rect 75460 347064 75512 347070
rect 75460 347006 75512 347012
rect 73252 346724 73304 346730
rect 73252 346666 73304 346672
rect 69296 346588 69348 346594
rect 69296 346530 69348 346536
rect 65984 346248 66036 346254
rect 65984 346190 66036 346196
rect 69308 344894 69336 346530
rect 75472 346497 75500 347006
rect 76760 346662 76788 347414
rect 78048 347002 78076 347647
rect 79152 347002 79180 347647
rect 81084 347206 81112 347647
rect 83660 347274 83688 347647
rect 83648 347268 83700 347274
rect 83648 347210 83700 347216
rect 81072 347200 81124 347206
rect 81072 347142 81124 347148
rect 78036 346996 78088 347002
rect 78036 346938 78088 346944
rect 79140 346996 79192 347002
rect 79140 346938 79192 346944
rect 76748 346656 76800 346662
rect 76748 346598 76800 346604
rect 79152 346526 79180 346938
rect 79140 346520 79192 346526
rect 75458 346488 75514 346497
rect 79140 346462 79192 346468
rect 75458 346423 75514 346432
rect 96080 346186 96108 347647
rect 100956 347138 100984 347647
rect 100944 347132 100996 347138
rect 100944 347074 100996 347080
rect 96068 346180 96120 346186
rect 96068 346122 96120 346128
rect 106108 346118 106136 347647
rect 106096 346112 106148 346118
rect 106096 346054 106148 346060
rect 108684 346050 108712 347647
rect 108672 346044 108724 346050
rect 108672 345986 108724 345992
rect 111076 345982 111104 347647
rect 111064 345976 111116 345982
rect 111064 345918 111116 345924
rect 113468 345846 113496 347647
rect 115860 345914 115888 347647
rect 115848 345908 115900 345914
rect 115848 345850 115900 345856
rect 113456 345840 113508 345846
rect 113456 345782 113508 345788
rect 118620 345778 118648 347647
rect 118608 345772 118660 345778
rect 118608 345714 118660 345720
rect 121012 345710 121040 347647
rect 123404 346866 123432 347647
rect 125980 346934 126008 347647
rect 125968 346928 126020 346934
rect 125968 346870 126020 346876
rect 123392 346860 123444 346866
rect 123392 346802 123444 346808
rect 121000 345704 121052 345710
rect 121000 345646 121052 345652
rect 69296 344888 69348 344894
rect 69296 344830 69348 344836
rect 150990 335472 151046 335481
rect 150990 335407 151046 335416
rect 151004 335374 151032 335407
rect 150992 335368 151044 335374
rect 150992 335310 151044 335316
rect 60832 334620 60884 334626
rect 60832 334562 60884 334568
rect 93490 249792 93546 249801
rect 93490 249727 93546 249736
rect 95882 249792 95938 249801
rect 95882 249727 95938 249736
rect 98550 249792 98606 249801
rect 98550 249727 98606 249736
rect 103518 249792 103574 249801
rect 103518 249727 103574 249736
rect 106002 249792 106058 249801
rect 106002 249727 106058 249736
rect 108578 249792 108634 249801
rect 108578 249727 108634 249736
rect 111062 249792 111118 249801
rect 111062 249727 111064 249736
rect 50802 249656 50858 249665
rect 50802 249591 50858 249600
rect 53654 249656 53710 249665
rect 53654 249591 53710 249600
rect 56046 249656 56102 249665
rect 56046 249591 56102 249600
rect 58530 249656 58586 249665
rect 58530 249591 58586 249600
rect 50816 249082 50844 249591
rect 53668 249150 53696 249591
rect 56060 249218 56088 249591
rect 58544 249286 58572 249591
rect 93504 249354 93532 249727
rect 95896 249422 95924 249727
rect 98564 249490 98592 249727
rect 103532 249558 103560 249727
rect 106016 249626 106044 249727
rect 108592 249694 108620 249727
rect 111116 249727 111118 249736
rect 111064 249698 111116 249704
rect 108580 249688 108632 249694
rect 108580 249630 108632 249636
rect 113454 249656 113510 249665
rect 106004 249620 106056 249626
rect 113454 249591 113510 249600
rect 115846 249656 115902 249665
rect 115846 249591 115902 249600
rect 120906 249656 120962 249665
rect 120906 249591 120962 249600
rect 106004 249562 106056 249568
rect 103520 249552 103572 249558
rect 103520 249494 103572 249500
rect 98552 249484 98604 249490
rect 98552 249426 98604 249432
rect 95884 249416 95936 249422
rect 95884 249358 95936 249364
rect 93492 249348 93544 249354
rect 93492 249290 93544 249296
rect 58532 249280 58584 249286
rect 58532 249222 58584 249228
rect 56048 249212 56100 249218
rect 56048 249154 56100 249160
rect 53656 249144 53708 249150
rect 53656 249086 53708 249092
rect 45928 249076 45980 249082
rect 45928 249018 45980 249024
rect 50804 249076 50856 249082
rect 50804 249018 50856 249024
rect 36452 248328 36504 248334
rect 35898 248296 35954 248305
rect 29552 248260 29604 248266
rect 35898 248231 35954 248240
rect 36450 248296 36452 248305
rect 36504 248296 36506 248305
rect 36450 248231 36506 248240
rect 38658 248296 38714 248305
rect 38658 248231 38660 248240
rect 29552 248202 29604 248208
rect 19984 248056 20036 248062
rect 19984 247998 20036 248004
rect 19892 247988 19944 247994
rect 19892 247930 19944 247936
rect 19800 247920 19852 247926
rect 19800 247862 19852 247868
rect 19708 148436 19760 148442
rect 19708 148378 19760 148384
rect 19708 147892 19760 147898
rect 19708 147834 19760 147840
rect 19720 147694 19748 147834
rect 19708 147688 19760 147694
rect 19708 147630 19760 147636
rect 19812 147286 19840 247862
rect 19904 147354 19932 247930
rect 19996 247110 20024 247998
rect 29564 247761 29592 248202
rect 35912 248198 35940 248231
rect 38712 248231 38714 248240
rect 44178 248296 44234 248305
rect 45940 248266 45968 249018
rect 113468 249014 113496 249591
rect 113456 249008 113508 249014
rect 113456 248950 113508 248956
rect 115860 248946 115888 249591
rect 115848 248940 115900 248946
rect 115848 248882 115900 248888
rect 120920 248878 120948 249591
rect 120908 248872 120960 248878
rect 120908 248814 120960 248820
rect 50160 248396 50212 248402
rect 50160 248338 50212 248344
rect 61200 248396 61252 248402
rect 61200 248338 61252 248344
rect 50172 248305 50200 248338
rect 61212 248305 61240 248338
rect 63592 248328 63644 248334
rect 46662 248296 46718 248305
rect 44178 248231 44234 248240
rect 45928 248260 45980 248266
rect 38660 248202 38712 248208
rect 44192 248198 44220 248231
rect 46662 248231 46664 248240
rect 45928 248202 45980 248208
rect 46716 248231 46718 248240
rect 50158 248296 50214 248305
rect 50158 248231 50214 248240
rect 61198 248296 61254 248305
rect 61198 248231 61254 248240
rect 61382 248296 61438 248305
rect 61382 248231 61438 248240
rect 62118 248296 62174 248305
rect 62118 248231 62174 248240
rect 63590 248296 63592 248305
rect 63644 248296 63646 248305
rect 63590 248231 63646 248240
rect 64878 248296 64934 248305
rect 64878 248231 64880 248240
rect 46664 248202 46716 248208
rect 35900 248192 35952 248198
rect 44180 248192 44232 248198
rect 35900 248134 35952 248140
rect 37278 248160 37334 248169
rect 40038 248160 40094 248169
rect 37278 248095 37280 248104
rect 37332 248095 37334 248104
rect 38108 248124 38160 248130
rect 37280 248066 37332 248072
rect 40038 248095 40094 248104
rect 41418 248160 41474 248169
rect 41418 248095 41420 248104
rect 38108 248066 38160 248072
rect 29550 247752 29606 247761
rect 29550 247687 29606 247696
rect 38120 247625 38148 248066
rect 40052 248062 40080 248095
rect 41472 248095 41474 248104
rect 43074 248160 43130 248169
rect 44180 248134 44232 248140
rect 45282 248160 45338 248169
rect 43074 248095 43130 248104
rect 41420 248066 41472 248072
rect 40040 248056 40092 248062
rect 40040 247998 40092 248004
rect 43088 247994 43116 248095
rect 43076 247988 43128 247994
rect 43076 247930 43128 247936
rect 44192 247926 44220 248134
rect 45282 248095 45338 248104
rect 47582 248160 47638 248169
rect 47582 248095 47638 248104
rect 45296 247994 45324 248095
rect 44272 247988 44324 247994
rect 44272 247930 44324 247936
rect 45284 247988 45336 247994
rect 45284 247930 45336 247936
rect 44180 247920 44232 247926
rect 44180 247862 44232 247868
rect 44284 247654 44312 247930
rect 47596 247858 47624 248095
rect 50172 247926 50200 248231
rect 59452 248124 59504 248130
rect 59452 248066 59504 248072
rect 50160 247920 50212 247926
rect 48686 247888 48742 247897
rect 47584 247852 47636 247858
rect 59464 247897 59492 248066
rect 61396 248062 61424 248231
rect 62132 248198 62160 248231
rect 64932 248231 64934 248240
rect 65982 248296 66038 248305
rect 65982 248231 66038 248240
rect 67638 248296 67694 248305
rect 67638 248231 67694 248240
rect 70950 248296 71006 248305
rect 70950 248231 71006 248240
rect 73802 248296 73858 248305
rect 73802 248231 73804 248240
rect 64880 248202 64932 248208
rect 65996 248198 66024 248231
rect 62120 248192 62172 248198
rect 62120 248134 62172 248140
rect 65984 248192 66036 248198
rect 65984 248134 66036 248140
rect 61384 248056 61436 248062
rect 61384 247998 61436 248004
rect 63498 248024 63554 248033
rect 63498 247959 63500 247968
rect 63552 247959 63554 247968
rect 63500 247930 63552 247936
rect 67652 247926 67680 248231
rect 68376 248056 68428 248062
rect 68376 247998 68428 248004
rect 67640 247920 67692 247926
rect 50160 247862 50212 247868
rect 58070 247888 58126 247897
rect 48686 247823 48742 247832
rect 58070 247823 58126 247832
rect 59450 247888 59506 247897
rect 59450 247823 59506 247832
rect 66258 247888 66314 247897
rect 68388 247897 68416 247998
rect 70964 247994 70992 248231
rect 73856 248231 73858 248240
rect 77298 248296 77354 248305
rect 77298 248231 77354 248240
rect 78494 248296 78550 248305
rect 78494 248231 78550 248240
rect 83646 248296 83702 248305
rect 83646 248231 83702 248240
rect 73804 248202 73856 248208
rect 77312 248130 77340 248231
rect 78508 248130 78536 248231
rect 77300 248124 77352 248130
rect 77300 248066 77352 248072
rect 78496 248124 78548 248130
rect 78496 248066 78548 248072
rect 81070 248024 81126 248033
rect 70952 247988 71004 247994
rect 81070 247959 81126 247968
rect 70952 247930 71004 247936
rect 67640 247862 67692 247868
rect 67730 247888 67786 247897
rect 66258 247823 66260 247832
rect 47584 247794 47636 247800
rect 48700 247790 48728 247823
rect 48688 247784 48740 247790
rect 48688 247726 48740 247732
rect 58084 247722 58112 247823
rect 58072 247716 58124 247722
rect 58072 247658 58124 247664
rect 44272 247648 44324 247654
rect 38106 247616 38162 247625
rect 44272 247590 44324 247596
rect 38106 247551 38162 247560
rect 52366 247480 52422 247489
rect 52422 247438 52592 247466
rect 59464 247450 59492 247823
rect 66312 247823 66314 247832
rect 67730 247823 67786 247832
rect 68374 247888 68430 247897
rect 68374 247823 68430 247832
rect 76102 247888 76158 247897
rect 76102 247823 76158 247832
rect 66260 247794 66312 247800
rect 67744 247790 67772 247823
rect 67732 247784 67784 247790
rect 67732 247726 67784 247732
rect 74998 247752 75054 247761
rect 74998 247687 75054 247696
rect 75918 247752 75974 247761
rect 75918 247687 75920 247696
rect 75012 247654 75040 247687
rect 75972 247687 75974 247696
rect 75920 247658 75972 247664
rect 76116 247654 76144 247823
rect 63224 247648 63276 247654
rect 75000 247648 75052 247654
rect 63224 247590 63276 247596
rect 71778 247616 71834 247625
rect 52366 247415 52422 247424
rect 52564 247382 52592 247438
rect 59452 247444 59504 247450
rect 59452 247386 59504 247392
rect 52552 247376 52604 247382
rect 52552 247318 52604 247324
rect 53746 247344 53802 247353
rect 52460 247308 52512 247314
rect 52460 247250 52512 247256
rect 19984 247104 20036 247110
rect 19984 247046 20036 247052
rect 52366 247072 52422 247081
rect 52472 247058 52500 247250
rect 52422 247030 52500 247058
rect 52366 247007 52422 247016
rect 52472 235754 52500 247030
rect 52460 235748 52512 235754
rect 52460 235690 52512 235696
rect 52564 235618 52592 247318
rect 53802 247302 53880 247330
rect 53746 247279 53802 247288
rect 53852 247246 53880 247302
rect 53840 247240 53892 247246
rect 53840 247182 53892 247188
rect 53852 235822 53880 247182
rect 55128 247172 55180 247178
rect 55128 247114 55180 247120
rect 55140 247081 55168 247114
rect 56612 247110 56640 247141
rect 56600 247104 56652 247110
rect 55126 247072 55182 247081
rect 56506 247072 56562 247081
rect 55182 247030 55260 247058
rect 55126 247007 55182 247016
rect 53840 235816 53892 235822
rect 53840 235758 53892 235764
rect 55232 235686 55260 247030
rect 56562 247052 56600 247058
rect 63236 247081 63264 247590
rect 75000 247590 75052 247596
rect 76104 247648 76156 247654
rect 76104 247590 76156 247596
rect 81084 247586 81112 247959
rect 83660 247926 83688 248231
rect 86038 248024 86094 248033
rect 86038 247959 86094 247968
rect 88246 248024 88302 248033
rect 88246 247959 88302 247968
rect 91006 248024 91062 248033
rect 91006 247959 91062 247968
rect 101218 248024 101274 248033
rect 101218 247959 101274 247968
rect 83648 247920 83700 247926
rect 83648 247862 83700 247868
rect 86052 247858 86080 247959
rect 86040 247852 86092 247858
rect 86040 247794 86092 247800
rect 88260 247790 88288 247959
rect 88248 247784 88300 247790
rect 88248 247726 88300 247732
rect 91020 247722 91048 247959
rect 91008 247716 91060 247722
rect 91008 247658 91060 247664
rect 71778 247551 71834 247560
rect 81072 247580 81124 247586
rect 69018 247480 69074 247489
rect 69018 247415 69074 247424
rect 69032 247382 69060 247415
rect 69020 247376 69072 247382
rect 69020 247318 69072 247324
rect 70398 247344 70454 247353
rect 70398 247279 70400 247288
rect 70452 247279 70454 247288
rect 70400 247250 70452 247256
rect 71792 247246 71820 247551
rect 81072 247522 81124 247528
rect 101232 247518 101260 247959
rect 101220 247512 101272 247518
rect 101220 247454 101272 247460
rect 73250 247344 73306 247353
rect 73250 247279 73306 247288
rect 71780 247240 71832 247246
rect 71780 247182 71832 247188
rect 73158 247208 73214 247217
rect 73158 247143 73160 247152
rect 73212 247143 73214 247152
rect 73160 247114 73212 247120
rect 73264 247110 73292 247279
rect 73252 247104 73304 247110
rect 56562 247046 56652 247052
rect 57978 247072 58034 247081
rect 56562 247030 56640 247046
rect 56506 247007 56562 247016
rect 56612 235890 56640 247030
rect 57978 247007 58034 247016
rect 63222 247072 63278 247081
rect 73252 247046 73304 247052
rect 63222 247007 63278 247016
rect 56600 235884 56652 235890
rect 56600 235826 56652 235832
rect 55220 235680 55272 235686
rect 55220 235622 55272 235628
rect 52552 235612 52604 235618
rect 52552 235554 52604 235560
rect 57992 235278 58020 247007
rect 150440 235952 150492 235958
rect 150440 235894 150492 235900
rect 57980 235272 58032 235278
rect 57980 235214 58032 235220
rect 150452 234705 150480 235894
rect 150438 234696 150494 234705
rect 150438 234631 150440 234640
rect 150492 234631 150494 234640
rect 150440 234602 150492 234608
rect 150452 234571 150480 234602
rect 48318 149560 48374 149569
rect 48318 149495 48374 149504
rect 50802 149560 50858 149569
rect 50802 149495 50858 149504
rect 56046 149560 56102 149569
rect 56046 149495 56102 149504
rect 58530 149560 58586 149569
rect 58530 149495 58586 149504
rect 60646 149560 60702 149569
rect 60646 149495 60702 149504
rect 71226 149560 71282 149569
rect 71226 149495 71282 149504
rect 73618 149560 73674 149569
rect 73618 149495 73674 149504
rect 83554 149560 83610 149569
rect 83554 149495 83610 149504
rect 93490 149560 93546 149569
rect 93490 149495 93546 149504
rect 98550 149560 98606 149569
rect 98550 149495 98606 149504
rect 103518 149560 103574 149569
rect 103518 149495 103574 149504
rect 113454 149560 113510 149569
rect 113454 149495 113510 149504
rect 115846 149560 115902 149569
rect 115846 149495 115902 149504
rect 120906 149560 120962 149569
rect 120906 149495 120962 149504
rect 19984 148436 20036 148442
rect 19984 148378 20036 148384
rect 19996 147898 20024 148378
rect 48332 148374 48360 149495
rect 50816 148442 50844 149495
rect 53654 149016 53710 149025
rect 53654 148951 53710 148960
rect 53668 148510 53696 148951
rect 56060 148578 56088 149495
rect 58544 148646 58572 149495
rect 60660 148714 60688 149495
rect 60648 148708 60700 148714
rect 60648 148650 60700 148656
rect 58532 148640 58584 148646
rect 58532 148582 58584 148588
rect 56048 148572 56100 148578
rect 56048 148514 56100 148520
rect 53656 148504 53708 148510
rect 53656 148446 53708 148452
rect 50804 148436 50856 148442
rect 50804 148378 50856 148384
rect 48320 148368 48372 148374
rect 48320 148310 48372 148316
rect 19984 147892 20036 147898
rect 19984 147834 20036 147840
rect 48228 147892 48280 147898
rect 48228 147834 48280 147840
rect 19892 147348 19944 147354
rect 19892 147290 19944 147296
rect 19800 147280 19852 147286
rect 19522 147248 19578 147257
rect 19800 147222 19852 147228
rect 19522 147183 19578 147192
rect 19536 147098 19564 147183
rect 19708 147144 19760 147150
rect 19536 147070 19656 147098
rect 19708 147086 19760 147092
rect 19444 142126 19564 142154
rect 19536 48113 19564 142126
rect 19628 48210 19656 147070
rect 19616 48204 19668 48210
rect 19616 48146 19668 48152
rect 19522 48104 19578 48113
rect 19522 48039 19578 48048
rect 19340 47728 19392 47734
rect 19340 47670 19392 47676
rect 18512 47534 18564 47540
rect 18970 47560 19026 47569
rect 18970 47495 19026 47504
rect 19720 47462 19748 147086
rect 19812 47530 19840 147222
rect 19904 147150 19932 147290
rect 19892 147144 19944 147150
rect 19892 147086 19944 147092
rect 19996 47802 20024 147834
rect 48136 147824 48188 147830
rect 48136 147766 48188 147772
rect 35898 147656 35954 147665
rect 35898 147591 35954 147600
rect 37002 147656 37058 147665
rect 37002 147591 37004 147600
rect 20628 147552 20680 147558
rect 20628 147494 20680 147500
rect 20640 146334 20668 147494
rect 35912 147490 35940 147591
rect 37056 147591 37058 147600
rect 38106 147656 38162 147665
rect 38106 147591 38162 147600
rect 39578 147656 39634 147665
rect 39578 147591 39634 147600
rect 43074 147656 43130 147665
rect 43074 147591 43130 147600
rect 44178 147656 44234 147665
rect 44178 147591 44234 147600
rect 45282 147656 45338 147665
rect 45282 147591 45338 147600
rect 46570 147656 46626 147665
rect 46570 147591 46626 147600
rect 47674 147656 47730 147665
rect 47674 147591 47730 147600
rect 37004 147562 37056 147568
rect 35900 147484 35952 147490
rect 35900 147426 35952 147432
rect 38120 147422 38148 147591
rect 38108 147416 38160 147422
rect 38108 147358 38160 147364
rect 21364 147144 21416 147150
rect 21364 147086 21416 147092
rect 21376 146946 21404 147086
rect 21364 146940 21416 146946
rect 21364 146882 21416 146888
rect 39592 146538 39620 147591
rect 43088 147354 43116 147591
rect 43076 147348 43128 147354
rect 43076 147290 43128 147296
rect 44192 147286 44220 147591
rect 44180 147280 44232 147286
rect 44180 147222 44232 147228
rect 44732 147280 44784 147286
rect 44732 147222 44784 147228
rect 44744 146674 44772 147222
rect 45296 146742 45324 147591
rect 46584 147286 46612 147591
rect 47688 147422 47716 147591
rect 48148 147490 48176 147766
rect 48240 147626 48268 147834
rect 58072 147756 58124 147762
rect 58072 147698 58124 147704
rect 59360 147756 59412 147762
rect 59360 147698 59412 147704
rect 58084 147665 58112 147698
rect 48686 147656 48742 147665
rect 48228 147620 48280 147626
rect 48686 147591 48742 147600
rect 50158 147656 50214 147665
rect 50158 147591 50160 147600
rect 48228 147562 48280 147568
rect 48136 147484 48188 147490
rect 48136 147426 48188 147432
rect 47676 147416 47728 147422
rect 47676 147358 47728 147364
rect 46020 147280 46072 147286
rect 46020 147222 46072 147228
rect 46572 147280 46624 147286
rect 46572 147222 46624 147228
rect 45284 146736 45336 146742
rect 45284 146678 45336 146684
rect 44732 146668 44784 146674
rect 44732 146610 44784 146616
rect 39580 146532 39632 146538
rect 39580 146474 39632 146480
rect 46032 146402 46060 147222
rect 46020 146396 46072 146402
rect 46020 146338 46072 146344
rect 47688 146334 47716 147358
rect 48700 147218 48728 147591
rect 50212 147591 50214 147600
rect 51446 147656 51502 147665
rect 51446 147591 51502 147600
rect 52274 147656 52330 147665
rect 52274 147591 52330 147600
rect 53378 147656 53434 147665
rect 53378 147591 53434 147600
rect 54022 147656 54078 147665
rect 54022 147591 54078 147600
rect 56046 147656 56102 147665
rect 56046 147591 56102 147600
rect 58070 147656 58126 147665
rect 58070 147591 58126 147600
rect 50160 147562 50212 147568
rect 48688 147212 48740 147218
rect 48688 147154 48740 147160
rect 50172 146878 50200 147562
rect 51460 147490 51488 147591
rect 51448 147484 51500 147490
rect 51448 147426 51500 147432
rect 50160 146872 50212 146878
rect 50160 146814 50212 146820
rect 51460 146810 51488 147426
rect 52288 147082 52316 147591
rect 52276 147076 52328 147082
rect 52276 147018 52328 147024
rect 53392 147014 53420 147591
rect 54036 147150 54064 147591
rect 54024 147144 54076 147150
rect 54024 147086 54076 147092
rect 53380 147008 53432 147014
rect 53380 146950 53432 146956
rect 51448 146804 51500 146810
rect 51448 146746 51500 146752
rect 54036 146606 54064 147086
rect 56060 146946 56088 147591
rect 59372 147354 59400 147698
rect 59556 147694 59584 147725
rect 59544 147688 59596 147694
rect 59542 147656 59544 147665
rect 59596 147656 59598 147665
rect 59542 147591 59598 147600
rect 59556 147490 59584 147591
rect 60660 147529 60688 148650
rect 61658 147656 61714 147665
rect 61658 147591 61714 147600
rect 62762 147656 62818 147665
rect 62762 147591 62818 147600
rect 63590 147656 63646 147665
rect 63590 147591 63592 147600
rect 61672 147558 61700 147591
rect 61660 147552 61712 147558
rect 60646 147520 60702 147529
rect 59544 147484 59596 147490
rect 61660 147494 61712 147500
rect 60646 147455 60702 147464
rect 59544 147426 59596 147432
rect 59360 147348 59412 147354
rect 59360 147290 59412 147296
rect 56048 146940 56100 146946
rect 56048 146882 56100 146888
rect 62776 146674 62804 147591
rect 63644 147591 63646 147600
rect 63866 147656 63922 147665
rect 63866 147591 63922 147600
rect 65154 147656 65210 147665
rect 65154 147591 65210 147600
rect 66166 147656 66222 147665
rect 66166 147591 66222 147600
rect 66350 147656 66406 147665
rect 66350 147591 66406 147600
rect 67638 147656 67694 147665
rect 67638 147591 67694 147600
rect 68282 147656 68338 147665
rect 68282 147591 68338 147600
rect 68466 147656 68522 147665
rect 68466 147591 68522 147600
rect 69754 147656 69810 147665
rect 69754 147591 69810 147600
rect 63592 147562 63644 147568
rect 63880 146742 63908 147591
rect 65168 147286 65196 147591
rect 66180 147558 66208 147591
rect 66168 147552 66220 147558
rect 66168 147494 66220 147500
rect 66364 147422 66392 147591
rect 66352 147416 66404 147422
rect 66352 147358 66404 147364
rect 65156 147280 65208 147286
rect 65156 147222 65208 147228
rect 67652 147218 67680 147591
rect 68296 147218 68324 147591
rect 67640 147212 67692 147218
rect 67640 147154 67692 147160
rect 68284 147212 68336 147218
rect 68284 147154 68336 147160
rect 68480 146878 68508 147591
rect 68468 146872 68520 146878
rect 68468 146814 68520 146820
rect 69768 146810 69796 147591
rect 70400 147416 70452 147422
rect 70400 147358 70452 147364
rect 70412 147257 70440 147358
rect 70398 147248 70454 147257
rect 70398 147183 70454 147192
rect 71042 147248 71098 147257
rect 71042 147183 71098 147192
rect 71056 147082 71084 147183
rect 71240 147150 71268 149495
rect 73632 148714 73660 149495
rect 76102 149016 76158 149025
rect 76102 148951 76158 148960
rect 76116 148782 76144 148951
rect 83568 148850 83596 149495
rect 86038 149016 86094 149025
rect 93504 148986 93532 149495
rect 98564 149054 98592 149495
rect 98552 149048 98604 149054
rect 98552 148990 98604 148996
rect 86038 148951 86094 148960
rect 93492 148980 93544 148986
rect 86052 148918 86080 148951
rect 93492 148922 93544 148928
rect 86040 148912 86092 148918
rect 86040 148854 86092 148860
rect 83556 148844 83608 148850
rect 83556 148786 83608 148792
rect 76104 148776 76156 148782
rect 76104 148718 76156 148724
rect 73620 148708 73672 148714
rect 73620 148650 73672 148656
rect 72146 147656 72202 147665
rect 72146 147591 72202 147600
rect 73250 147656 73306 147665
rect 73250 147591 73306 147600
rect 73710 147656 73766 147665
rect 73710 147591 73766 147600
rect 75642 147656 75698 147665
rect 75642 147591 75698 147600
rect 76930 147656 76986 147665
rect 76930 147591 76986 147600
rect 78034 147656 78090 147665
rect 78034 147591 78090 147600
rect 78494 147656 78550 147665
rect 78494 147591 78550 147600
rect 79138 147656 79194 147665
rect 79138 147591 79194 147600
rect 81070 147656 81126 147665
rect 81070 147591 81126 147600
rect 88246 147656 88302 147665
rect 88246 147591 88302 147600
rect 91006 147656 91062 147665
rect 91006 147591 91062 147600
rect 95974 147656 96030 147665
rect 95974 147591 96030 147600
rect 100942 147656 100998 147665
rect 100942 147591 100998 147600
rect 71228 147144 71280 147150
rect 71228 147086 71280 147092
rect 71044 147076 71096 147082
rect 71044 147018 71096 147024
rect 72160 147014 72188 147591
rect 72148 147008 72200 147014
rect 72148 146950 72200 146956
rect 69756 146804 69808 146810
rect 69756 146746 69808 146752
rect 63868 146736 63920 146742
rect 63868 146678 63920 146684
rect 62764 146668 62816 146674
rect 62764 146610 62816 146616
rect 73264 146606 73292 147591
rect 73724 146946 73752 147591
rect 75656 147422 75684 147591
rect 75826 147520 75882 147529
rect 75826 147455 75882 147464
rect 75840 147422 75868 147455
rect 75644 147416 75696 147422
rect 75644 147358 75696 147364
rect 75828 147416 75880 147422
rect 75828 147358 75880 147364
rect 76944 147354 76972 147591
rect 78048 147490 78076 147591
rect 78508 147490 78536 147591
rect 78036 147484 78088 147490
rect 78036 147426 78088 147432
rect 78496 147484 78548 147490
rect 78496 147426 78548 147432
rect 79152 147422 79180 147591
rect 81084 147422 81112 147591
rect 79140 147416 79192 147422
rect 79140 147358 79192 147364
rect 81072 147416 81124 147422
rect 81072 147358 81124 147364
rect 88260 147354 88288 147591
rect 76932 147348 76984 147354
rect 76932 147290 76984 147296
rect 88248 147348 88300 147354
rect 88248 147290 88300 147296
rect 91020 147286 91048 147591
rect 91008 147280 91060 147286
rect 91008 147222 91060 147228
rect 95988 147082 96016 147591
rect 95976 147076 96028 147082
rect 95976 147018 96028 147024
rect 100956 146946 100984 147591
rect 103532 147014 103560 149495
rect 113468 148306 113496 149495
rect 113456 148300 113508 148306
rect 113456 148242 113508 148248
rect 115860 148238 115888 149495
rect 115848 148232 115900 148238
rect 115848 148174 115900 148180
rect 120920 148170 120948 149495
rect 120908 148164 120960 148170
rect 120908 148106 120960 148112
rect 106094 147656 106150 147665
rect 106094 147591 106150 147600
rect 108854 147656 108910 147665
rect 108854 147591 108910 147600
rect 111614 147656 111670 147665
rect 111614 147591 111670 147600
rect 103520 147008 103572 147014
rect 103520 146950 103572 146956
rect 73712 146940 73764 146946
rect 73712 146882 73764 146888
rect 100944 146940 100996 146946
rect 100944 146882 100996 146888
rect 106108 146878 106136 147591
rect 106096 146872 106148 146878
rect 106096 146814 106148 146820
rect 108868 146810 108896 147591
rect 108856 146804 108908 146810
rect 108856 146746 108908 146752
rect 111628 146742 111656 147591
rect 156616 146878 156644 450055
rect 156708 346866 156736 459614
rect 157982 456376 158038 456385
rect 157982 456311 158038 456320
rect 157890 452296 157946 452305
rect 156972 452260 157024 452266
rect 157890 452231 157946 452240
rect 156972 452202 157024 452208
rect 156880 451444 156932 451450
rect 156880 451386 156932 451392
rect 156786 450528 156842 450537
rect 156786 450463 156842 450472
rect 156696 346860 156748 346866
rect 156696 346802 156748 346808
rect 156696 235952 156748 235958
rect 156696 235894 156748 235900
rect 156708 234666 156736 235894
rect 156696 234660 156748 234666
rect 156696 234602 156748 234608
rect 156604 146872 156656 146878
rect 156604 146814 156656 146820
rect 111616 146736 111668 146742
rect 111616 146678 111668 146684
rect 54024 146600 54076 146606
rect 54024 146542 54076 146548
rect 73252 146600 73304 146606
rect 73252 146542 73304 146548
rect 20628 146328 20680 146334
rect 20628 146270 20680 146276
rect 47676 146328 47728 146334
rect 47676 146270 47728 146276
rect 156708 136610 156736 234602
rect 156800 147529 156828 450463
rect 156892 348974 156920 451386
rect 156880 348968 156932 348974
rect 156880 348910 156932 348916
rect 156984 348906 157012 452202
rect 157800 451784 157852 451790
rect 157800 451726 157852 451732
rect 157812 349110 157840 451726
rect 157800 349104 157852 349110
rect 157800 349046 157852 349052
rect 156972 348900 157024 348906
rect 156972 348842 157024 348848
rect 157904 348294 157932 452231
rect 157892 348288 157944 348294
rect 157892 348230 157944 348236
rect 156786 147520 156842 147529
rect 156786 147455 156842 147464
rect 157996 146742 158024 456311
rect 158076 455796 158128 455802
rect 158076 455738 158128 455744
rect 158088 247586 158116 455738
rect 158260 455728 158312 455734
rect 158260 455670 158312 455676
rect 158166 455560 158222 455569
rect 158166 455495 158222 455504
rect 158076 247580 158128 247586
rect 158076 247522 158128 247528
rect 158180 146810 158208 455495
rect 158272 247654 158300 455670
rect 158628 451716 158680 451722
rect 158628 451658 158680 451664
rect 158534 451616 158590 451625
rect 158534 451551 158590 451560
rect 158352 451512 158404 451518
rect 158352 451454 158404 451460
rect 158364 348634 158392 451454
rect 158444 451376 158496 451382
rect 158444 451318 158496 451324
rect 158352 348628 158404 348634
rect 158352 348570 158404 348576
rect 158456 348226 158484 451318
rect 158548 349042 158576 451551
rect 158536 349036 158588 349042
rect 158536 348978 158588 348984
rect 158640 348702 158668 451658
rect 158720 435396 158772 435402
rect 158720 435338 158772 435344
rect 158628 348696 158680 348702
rect 158628 348638 158680 348644
rect 158444 348220 158496 348226
rect 158444 348162 158496 348168
rect 158732 335306 158760 435338
rect 158810 429312 158866 429321
rect 158810 429247 158866 429256
rect 158720 335300 158772 335306
rect 158720 335242 158772 335248
rect 158732 334098 158760 335242
rect 158640 334070 158760 334098
rect 158260 247648 158312 247654
rect 158260 247590 158312 247596
rect 158640 235958 158668 334070
rect 158824 329769 158852 429247
rect 158810 329760 158866 329769
rect 158810 329695 158866 329704
rect 158824 316034 158852 329695
rect 158732 316006 158852 316034
rect 158628 235952 158680 235958
rect 158628 235894 158680 235900
rect 158732 230450 158760 316006
rect 158720 230444 158772 230450
rect 158720 230386 158772 230392
rect 158732 229265 158760 230386
rect 158718 229256 158774 229265
rect 158718 229191 158774 229200
rect 158168 146804 158220 146810
rect 158168 146746 158220 146752
rect 157984 146736 158036 146742
rect 157984 146678 158036 146684
rect 151268 136604 151320 136610
rect 151268 136546 151320 136552
rect 156696 136604 156748 136610
rect 156696 136546 156748 136552
rect 151280 135833 151308 136546
rect 151266 135824 151322 135833
rect 151266 135759 151322 135768
rect 158732 129713 158760 229191
rect 158718 129704 158774 129713
rect 158718 129639 158774 129648
rect 53472 49904 53524 49910
rect 53470 49872 53472 49881
rect 53524 49872 53526 49881
rect 60646 49872 60702 49881
rect 53470 49807 53526 49816
rect 59544 49836 59596 49842
rect 48318 49600 48374 49609
rect 48318 49535 48374 49544
rect 50802 49600 50858 49609
rect 50802 49535 50858 49544
rect 48332 49026 48360 49535
rect 50816 49094 50844 49535
rect 50804 49088 50856 49094
rect 50804 49030 50856 49036
rect 48320 49020 48372 49026
rect 48320 48962 48372 48968
rect 36820 48272 36872 48278
rect 36818 48240 36820 48249
rect 36872 48240 36874 48249
rect 36818 48175 36874 48184
rect 43166 48240 43222 48249
rect 43166 48175 43222 48184
rect 44178 48240 44234 48249
rect 44178 48175 44234 48184
rect 45374 48240 45430 48249
rect 45374 48175 45430 48184
rect 46570 48240 46626 48249
rect 46570 48175 46626 48184
rect 47582 48240 47638 48249
rect 47582 48175 47638 48184
rect 48686 48240 48742 48249
rect 48686 48175 48742 48184
rect 49698 48240 49754 48249
rect 49698 48175 49754 48184
rect 50250 48240 50306 48249
rect 50250 48175 50306 48184
rect 51446 48240 51502 48249
rect 51446 48175 51502 48184
rect 52366 48240 52422 48249
rect 52366 48175 52422 48184
rect 19984 47796 20036 47802
rect 19984 47738 20036 47744
rect 19800 47524 19852 47530
rect 19800 47466 19852 47472
rect 43180 47462 43208 48175
rect 44192 47530 44220 48175
rect 45388 47598 45416 48175
rect 46584 47666 46612 48175
rect 47596 47734 47624 48175
rect 48700 47938 48728 48175
rect 48688 47932 48740 47938
rect 48688 47874 48740 47880
rect 49712 47802 49740 48175
rect 49700 47796 49752 47802
rect 49700 47738 49752 47744
rect 47584 47728 47636 47734
rect 47584 47670 47636 47676
rect 48228 47728 48280 47734
rect 48228 47670 48280 47676
rect 46572 47660 46624 47666
rect 46572 47602 46624 47608
rect 48240 47598 48268 47670
rect 45376 47592 45428 47598
rect 45376 47534 45428 47540
rect 48228 47592 48280 47598
rect 48228 47534 48280 47540
rect 44180 47524 44232 47530
rect 44180 47466 44232 47472
rect 19708 47456 19760 47462
rect 19708 47398 19760 47404
rect 43168 47456 43220 47462
rect 43168 47398 43220 47404
rect 44192 47394 44220 47466
rect 44180 47388 44232 47394
rect 44180 47330 44232 47336
rect 18236 47320 18288 47326
rect 18236 47262 18288 47268
rect 50264 47258 50292 48175
rect 51460 47870 51488 48175
rect 51448 47864 51500 47870
rect 51448 47806 51500 47812
rect 50252 47252 50304 47258
rect 50252 47194 50304 47200
rect 51460 47122 51488 47806
rect 52380 47802 52408 48175
rect 53484 48006 53512 49807
rect 60646 49807 60702 49816
rect 59544 49778 59596 49784
rect 53654 49600 53710 49609
rect 53654 49535 53710 49544
rect 56046 49600 56102 49609
rect 56046 49535 56102 49544
rect 58530 49600 58586 49609
rect 58530 49535 58586 49544
rect 53668 49162 53696 49535
rect 56060 49230 56088 49535
rect 58544 49298 58572 49535
rect 58532 49292 58584 49298
rect 58532 49234 58584 49240
rect 56048 49224 56100 49230
rect 56048 49166 56100 49172
rect 53656 49156 53708 49162
rect 53656 49098 53708 49104
rect 59556 48278 59584 49778
rect 60660 49774 60688 49807
rect 60648 49768 60700 49774
rect 60648 49710 60700 49716
rect 91006 49736 91062 49745
rect 59544 48272 59596 48278
rect 54574 48240 54630 48249
rect 54574 48175 54630 48184
rect 55862 48240 55918 48249
rect 57978 48240 58034 48249
rect 55862 48175 55918 48184
rect 57060 48204 57112 48210
rect 53472 48000 53524 48006
rect 53472 47942 53524 47948
rect 54588 47938 54616 48175
rect 55876 48142 55904 48175
rect 57978 48175 58034 48184
rect 59542 48240 59544 48249
rect 59596 48240 59598 48249
rect 59542 48175 59598 48184
rect 57060 48146 57112 48152
rect 55864 48136 55916 48142
rect 55864 48078 55916 48084
rect 56508 48136 56560 48142
rect 56508 48078 56560 48084
rect 54576 47932 54628 47938
rect 54576 47874 54628 47880
rect 52368 47796 52420 47802
rect 52368 47738 52420 47744
rect 56520 47190 56548 48078
rect 57072 47569 57100 48146
rect 57058 47560 57114 47569
rect 57058 47495 57114 47504
rect 57992 47326 58020 48175
rect 60660 47977 60688 49710
rect 91006 49671 91062 49680
rect 95882 49736 95938 49745
rect 95882 49671 95884 49680
rect 91020 49638 91048 49671
rect 95936 49671 95938 49680
rect 95884 49642 95936 49648
rect 91008 49632 91060 49638
rect 80978 49600 81034 49609
rect 80978 49535 81034 49544
rect 83554 49600 83610 49609
rect 83554 49535 83610 49544
rect 86038 49600 86094 49609
rect 86038 49535 86094 49544
rect 88246 49600 88302 49609
rect 91008 49574 91060 49580
rect 98550 49600 98606 49609
rect 88246 49535 88248 49544
rect 80992 49366 81020 49535
rect 83568 49434 83596 49535
rect 86052 49502 86080 49535
rect 88300 49535 88302 49544
rect 98550 49535 98606 49544
rect 103518 49600 103574 49609
rect 103518 49535 103574 49544
rect 106002 49600 106058 49609
rect 106002 49535 106058 49544
rect 88248 49506 88300 49512
rect 86040 49496 86092 49502
rect 86040 49438 86092 49444
rect 83556 49428 83608 49434
rect 83556 49370 83608 49376
rect 80980 49360 81032 49366
rect 80980 49302 81032 49308
rect 98564 48958 98592 49535
rect 98552 48952 98604 48958
rect 98552 48894 98604 48900
rect 103532 48890 103560 49535
rect 103520 48884 103572 48890
rect 103520 48826 103572 48832
rect 106016 48822 106044 49535
rect 106004 48816 106056 48822
rect 106004 48758 106056 48764
rect 78036 48272 78088 48278
rect 61198 48240 61254 48249
rect 61198 48175 61200 48184
rect 61252 48175 61254 48184
rect 61382 48240 61438 48249
rect 61382 48175 61438 48184
rect 62210 48240 62266 48249
rect 62210 48175 62266 48184
rect 63958 48240 64014 48249
rect 63958 48175 64014 48184
rect 65062 48240 65118 48249
rect 65062 48175 65118 48184
rect 65982 48240 66038 48249
rect 65982 48175 66038 48184
rect 66258 48240 66314 48249
rect 66258 48175 66314 48184
rect 67638 48240 67694 48249
rect 67638 48175 67694 48184
rect 68374 48240 68430 48249
rect 68374 48175 68430 48184
rect 68558 48240 68614 48249
rect 68558 48175 68614 48184
rect 69754 48240 69810 48249
rect 69754 48175 69810 48184
rect 71134 48240 71190 48249
rect 71134 48175 71190 48184
rect 71778 48240 71834 48249
rect 71778 48175 71834 48184
rect 73250 48240 73306 48249
rect 73250 48175 73306 48184
rect 73802 48240 73858 48249
rect 73802 48175 73858 48184
rect 74354 48240 74410 48249
rect 74354 48175 74410 48184
rect 76102 48240 76158 48249
rect 76102 48175 76158 48184
rect 76378 48240 76434 48249
rect 76378 48175 76434 48184
rect 78034 48240 78036 48249
rect 125968 48272 126020 48278
rect 78088 48240 78090 48249
rect 78034 48175 78090 48184
rect 78494 48240 78550 48249
rect 78494 48175 78550 48184
rect 93582 48240 93638 48249
rect 93582 48175 93638 48184
rect 100942 48240 100998 48249
rect 100942 48175 100998 48184
rect 108854 48240 108910 48249
rect 108854 48175 108910 48184
rect 111154 48240 111210 48249
rect 111154 48175 111210 48184
rect 115846 48240 115902 48249
rect 115846 48175 115902 48184
rect 118606 48240 118662 48249
rect 118606 48175 118662 48184
rect 125966 48240 125968 48249
rect 126020 48240 126022 48249
rect 159376 48210 159404 463014
rect 159548 462936 159600 462942
rect 159548 462878 159600 462884
rect 159456 462800 159508 462806
rect 159456 462742 159508 462748
rect 125966 48175 126022 48184
rect 159364 48204 159416 48210
rect 61200 48146 61252 48152
rect 60646 47968 60702 47977
rect 60646 47903 60702 47912
rect 61396 47462 61424 48175
rect 61384 47456 61436 47462
rect 61384 47398 61436 47404
rect 62224 47394 62252 48175
rect 63866 48104 63922 48113
rect 63972 48074 64000 48175
rect 63866 48039 63922 48048
rect 63960 48068 64012 48074
rect 63880 47530 63908 48039
rect 63960 48010 64012 48016
rect 65076 47666 65104 48175
rect 65996 48142 66024 48175
rect 65984 48136 66036 48142
rect 65984 48078 66036 48084
rect 65064 47660 65116 47666
rect 65064 47602 65116 47608
rect 66272 47598 66300 48175
rect 67652 47734 67680 48175
rect 68388 47870 68416 48175
rect 68376 47864 68428 47870
rect 68376 47806 68428 47812
rect 67640 47728 67692 47734
rect 67640 47670 67692 47676
rect 66260 47592 66312 47598
rect 66260 47534 66312 47540
rect 63868 47524 63920 47530
rect 63868 47466 63920 47472
rect 62212 47388 62264 47394
rect 62212 47330 62264 47336
rect 57980 47320 58032 47326
rect 57980 47262 58032 47268
rect 68572 47258 68600 48175
rect 68560 47252 68612 47258
rect 68560 47194 68612 47200
rect 56508 47184 56560 47190
rect 56508 47126 56560 47132
rect 69768 47122 69796 48175
rect 71042 48104 71098 48113
rect 71042 48039 71098 48048
rect 71056 47802 71084 48039
rect 71148 47802 71176 48175
rect 71792 48006 71820 48175
rect 71780 48000 71832 48006
rect 71780 47942 71832 47948
rect 73264 47938 73292 48175
rect 73816 48006 73844 48175
rect 73804 48000 73856 48006
rect 73804 47942 73856 47948
rect 73252 47932 73304 47938
rect 73252 47874 73304 47880
rect 71044 47796 71096 47802
rect 71044 47738 71096 47744
rect 71136 47796 71188 47802
rect 71136 47738 71188 47744
rect 74368 47190 74396 48175
rect 76116 47938 76144 48175
rect 76104 47932 76156 47938
rect 76104 47874 76156 47880
rect 76392 47326 76420 48175
rect 78508 47734 78536 48175
rect 78496 47728 78548 47734
rect 78496 47670 78548 47676
rect 93596 47666 93624 48175
rect 93584 47660 93636 47666
rect 93584 47602 93636 47608
rect 100956 47598 100984 48175
rect 100944 47592 100996 47598
rect 100944 47534 100996 47540
rect 76380 47320 76432 47326
rect 76380 47262 76432 47268
rect 74356 47184 74408 47190
rect 74356 47126 74408 47132
rect 51448 47116 51500 47122
rect 51448 47058 51500 47064
rect 69756 47116 69808 47122
rect 69756 47058 69808 47064
rect 108868 46918 108896 48175
rect 111168 47530 111196 48175
rect 111156 47524 111208 47530
rect 111156 47466 111208 47472
rect 115860 47462 115888 48175
rect 115848 47456 115900 47462
rect 115848 47398 115900 47404
rect 118620 47394 118648 48175
rect 159364 48146 159416 48152
rect 159468 47870 159496 462742
rect 159560 48074 159588 462878
rect 159652 49298 159680 463082
rect 159640 49292 159692 49298
rect 159640 49234 159692 49240
rect 159744 49230 159772 463150
rect 159824 459740 159876 459746
rect 159824 459682 159876 459688
rect 159836 346934 159864 459682
rect 159824 346928 159876 346934
rect 159824 346870 159876 346876
rect 159732 49224 159784 49230
rect 159732 49166 159784 49172
rect 159548 48068 159600 48074
rect 159548 48010 159600 48016
rect 159456 47864 159508 47870
rect 159456 47806 159508 47812
rect 160756 47530 160784 465462
rect 161020 465452 161072 465458
rect 161020 465394 161072 465400
rect 160928 465384 160980 465390
rect 160928 465326 160980 465332
rect 160836 465316 160888 465322
rect 160836 465258 160888 465264
rect 160744 47524 160796 47530
rect 160744 47466 160796 47472
rect 160848 47394 160876 465258
rect 160940 47462 160968 465326
rect 161032 49473 161060 465394
rect 169024 464636 169076 464642
rect 169024 464578 169076 464584
rect 166724 464228 166776 464234
rect 166724 464170 166776 464176
rect 166356 464160 166408 464166
rect 166356 464102 166408 464108
rect 166630 464128 166686 464137
rect 163594 463992 163650 464001
rect 163594 463927 163650 463936
rect 162124 462732 162176 462738
rect 162124 462674 162176 462680
rect 161112 462664 161164 462670
rect 161112 462606 161164 462612
rect 161018 49464 161074 49473
rect 161018 49399 161074 49408
rect 161124 48142 161152 462606
rect 161204 461780 161256 461786
rect 161204 461722 161256 461728
rect 161216 49162 161244 461722
rect 161296 454504 161348 454510
rect 161296 454446 161348 454452
rect 161308 349586 161336 454446
rect 161296 349580 161348 349586
rect 161296 349522 161348 349528
rect 161480 89004 161532 89010
rect 161480 88946 161532 88952
rect 161204 49156 161256 49162
rect 161204 49098 161256 49104
rect 161112 48136 161164 48142
rect 161112 48078 161164 48084
rect 160928 47456 160980 47462
rect 160928 47398 160980 47404
rect 118608 47388 118660 47394
rect 118608 47330 118660 47336
rect 160836 47388 160888 47394
rect 160836 47330 160888 47336
rect 108856 46912 108908 46918
rect 108856 46854 108908 46860
rect 133880 46232 133932 46238
rect 133880 46174 133932 46180
rect 126980 42084 127032 42090
rect 126980 42026 127032 42032
rect 125600 39364 125652 39370
rect 125600 39306 125652 39312
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 1688 480 1716 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 39306
rect 126992 480 127020 42026
rect 130568 7608 130620 7614
rect 130568 7550 130620 7556
rect 128176 4820 128228 4826
rect 128176 4762 128228 4768
rect 128188 480 128216 4762
rect 130580 480 130608 7550
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 46174
rect 161492 16574 161520 88946
rect 162136 47802 162164 462674
rect 163502 462360 163558 462369
rect 163502 462295 163558 462304
rect 162492 459196 162544 459202
rect 162492 459138 162544 459144
rect 162400 457836 162452 457842
rect 162400 457778 162452 457784
rect 162308 456816 162360 456822
rect 162308 456758 162360 456764
rect 162216 455592 162268 455598
rect 162216 455534 162268 455540
rect 162228 147218 162256 455534
rect 162320 346050 162348 456758
rect 162412 346118 162440 457778
rect 162504 347070 162532 459138
rect 162768 457768 162820 457774
rect 162768 457710 162820 457716
rect 162676 456612 162728 456618
rect 162676 456554 162728 456560
rect 162584 456408 162636 456414
rect 162584 456350 162636 456356
rect 162492 347064 162544 347070
rect 162492 347006 162544 347012
rect 162400 346112 162452 346118
rect 162400 346054 162452 346060
rect 162308 346044 162360 346050
rect 162308 345986 162360 345992
rect 162596 345982 162624 456350
rect 162584 345976 162636 345982
rect 162584 345918 162636 345924
rect 162688 345846 162716 456554
rect 162780 349654 162808 457710
rect 163412 452192 163464 452198
rect 163412 452134 163464 452140
rect 162768 349648 162820 349654
rect 162768 349590 162820 349596
rect 163424 349382 163452 452134
rect 163412 349376 163464 349382
rect 163412 349318 163464 349324
rect 162676 345840 162728 345846
rect 162676 345782 162728 345788
rect 162216 147212 162268 147218
rect 162216 147154 162268 147160
rect 162124 47796 162176 47802
rect 162124 47738 162176 47744
rect 163516 46918 163544 462295
rect 163608 47598 163636 463927
rect 166264 463888 166316 463894
rect 163962 463856 164018 463865
rect 166264 463830 166316 463836
rect 163962 463791 164018 463800
rect 163778 463720 163834 463729
rect 163778 463655 163834 463664
rect 163688 462528 163740 462534
rect 163688 462470 163740 462476
rect 163700 48958 163728 462470
rect 163688 48952 163740 48958
rect 163688 48894 163740 48900
rect 163792 48822 163820 463655
rect 163870 456104 163926 456113
rect 163870 456039 163926 456048
rect 163884 49094 163912 456039
rect 163872 49088 163924 49094
rect 163872 49030 163924 49036
rect 163976 48890 164004 463791
rect 164148 460012 164200 460018
rect 164148 459954 164200 459960
rect 164056 455932 164108 455938
rect 164056 455874 164108 455880
rect 164068 147150 164096 455874
rect 164160 347002 164188 459954
rect 165160 456476 165212 456482
rect 165160 456418 165212 456424
rect 165068 456068 165120 456074
rect 165068 456010 165120 456016
rect 164976 455524 165028 455530
rect 164976 455466 165028 455472
rect 164884 455456 164936 455462
rect 164884 455398 164936 455404
rect 164148 346996 164200 347002
rect 164148 346938 164200 346944
rect 164896 345710 164924 455398
rect 164988 345778 165016 455466
rect 165080 346254 165108 456010
rect 165068 346248 165120 346254
rect 165068 346190 165120 346196
rect 165172 345914 165200 456418
rect 166172 451104 166224 451110
rect 166172 451046 166224 451052
rect 165252 450084 165304 450090
rect 165252 450026 165304 450032
rect 165160 345908 165212 345914
rect 165160 345850 165212 345856
rect 164976 345772 165028 345778
rect 164976 345714 165028 345720
rect 164884 345704 164936 345710
rect 164884 345646 164936 345652
rect 165264 344962 165292 450026
rect 165344 449608 165396 449614
rect 165344 449550 165396 449556
rect 165356 346322 165384 449550
rect 165344 346316 165396 346322
rect 165344 346258 165396 346264
rect 166184 346186 166212 451046
rect 166172 346180 166224 346186
rect 166172 346122 166224 346128
rect 165252 344956 165304 344962
rect 165252 344898 165304 344904
rect 165620 244996 165672 245002
rect 165620 244938 165672 244944
rect 164056 147144 164108 147150
rect 164056 147086 164108 147092
rect 163964 48884 164016 48890
rect 163964 48826 164016 48832
rect 163780 48816 163832 48822
rect 163780 48758 163832 48764
rect 163596 47592 163648 47598
rect 163596 47534 163648 47540
rect 163504 46912 163556 46918
rect 163504 46854 163556 46860
rect 165632 16574 165660 244938
rect 166276 47666 166304 463830
rect 166368 49434 166396 464102
rect 166630 464063 166686 464072
rect 166540 464024 166592 464030
rect 166540 463966 166592 463972
rect 166448 463956 166500 463962
rect 166448 463898 166500 463904
rect 166460 49638 166488 463898
rect 166448 49632 166500 49638
rect 166448 49574 166500 49580
rect 166552 49570 166580 463966
rect 166644 49706 166672 464063
rect 166632 49700 166684 49706
rect 166632 49642 166684 49648
rect 166540 49564 166592 49570
rect 166540 49506 166592 49512
rect 166356 49428 166408 49434
rect 166356 49370 166408 49376
rect 166736 49366 166764 464170
rect 166816 464092 166868 464098
rect 166816 464034 166868 464040
rect 166828 49502 166856 464034
rect 167736 463004 167788 463010
rect 167736 462946 167788 462952
rect 167644 456272 167696 456278
rect 167644 456214 167696 456220
rect 166908 454912 166960 454918
rect 166908 454854 166960 454860
rect 166920 348770 166948 454854
rect 166908 348764 166960 348770
rect 166908 348706 166960 348712
rect 166816 49496 166868 49502
rect 166816 49438 166868 49444
rect 166724 49360 166776 49366
rect 166724 49302 166776 49308
rect 166264 47660 166316 47666
rect 166264 47602 166316 47608
rect 167656 33114 167684 456214
rect 167748 45558 167776 462946
rect 167920 461916 167972 461922
rect 167920 461858 167972 461864
rect 167828 460488 167880 460494
rect 167828 460430 167880 460436
rect 167840 137970 167868 460430
rect 167932 241466 167960 461858
rect 168010 454744 168066 454753
rect 168010 454679 168066 454688
rect 168104 454708 168156 454714
rect 168024 344350 168052 454679
rect 168104 454650 168156 454656
rect 168116 344894 168144 454650
rect 168196 450696 168248 450702
rect 168196 450638 168248 450644
rect 168208 345030 168236 450638
rect 168196 345024 168248 345030
rect 168196 344966 168248 344972
rect 168104 344888 168156 344894
rect 168104 344830 168156 344836
rect 168012 344344 168064 344350
rect 168012 344286 168064 344292
rect 167920 241460 167972 241466
rect 167920 241402 167972 241408
rect 167828 137964 167880 137970
rect 167828 137906 167880 137912
rect 169036 47734 169064 464578
rect 171784 463820 171836 463826
rect 171784 463762 171836 463768
rect 170402 461544 170458 461553
rect 170402 461479 170458 461488
rect 169300 460556 169352 460562
rect 169300 460498 169352 460504
rect 169114 460184 169170 460193
rect 169114 460119 169170 460128
rect 169128 48006 169156 460119
rect 169206 458824 169262 458833
rect 169206 458759 169262 458768
rect 169116 48000 169168 48006
rect 169116 47942 169168 47948
rect 169220 47938 169248 458759
rect 169312 49026 169340 460498
rect 169392 456952 169444 456958
rect 169392 456894 169444 456900
rect 169404 247994 169432 456894
rect 169484 454776 169536 454782
rect 169484 454718 169536 454724
rect 169496 248198 169524 454718
rect 169668 454572 169720 454578
rect 169668 454514 169720 454520
rect 169574 452976 169630 452985
rect 169574 452911 169630 452920
rect 169484 248192 169536 248198
rect 169484 248134 169536 248140
rect 169588 248062 169616 452911
rect 169680 349518 169708 454514
rect 169668 349512 169720 349518
rect 169668 349454 169720 349460
rect 169576 248056 169628 248062
rect 169576 247998 169628 248004
rect 169392 247988 169444 247994
rect 169392 247930 169444 247936
rect 169300 49020 169352 49026
rect 169300 48962 169352 48968
rect 169208 47932 169260 47938
rect 169208 47874 169260 47880
rect 169024 47728 169076 47734
rect 169024 47670 169076 47676
rect 167736 45552 167788 45558
rect 167736 45494 167788 45500
rect 167644 33108 167696 33114
rect 167644 33050 167696 33056
rect 161492 16546 162072 16574
rect 165632 16546 166120 16574
rect 158904 3868 158956 3874
rect 158904 3810 158956 3816
rect 155408 3800 155460 3806
rect 155408 3742 155460 3748
rect 151820 3732 151872 3738
rect 151820 3674 151872 3680
rect 148324 3664 148376 3670
rect 148324 3606 148376 3612
rect 144736 3596 144788 3602
rect 144736 3538 144788 3544
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 137652 3460 137704 3466
rect 137652 3402 137704 3408
rect 137664 480 137692 3402
rect 141252 480 141280 3470
rect 144748 480 144776 3538
rect 148336 480 148364 3606
rect 151832 480 151860 3674
rect 155420 480 155448 3742
rect 158916 480 158944 3810
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 166092 480 166120 16546
rect 169576 8968 169628 8974
rect 169576 8910 169628 8916
rect 169588 480 169616 8910
rect 170416 6866 170444 461479
rect 170496 457496 170548 457502
rect 170496 457438 170548 457444
rect 170508 20670 170536 457438
rect 171796 247897 171824 463762
rect 174636 463344 174688 463350
rect 174636 463286 174688 463292
rect 174544 462596 174596 462602
rect 174544 462538 174596 462544
rect 172060 460420 172112 460426
rect 172060 460362 172112 460368
rect 171968 460352 172020 460358
rect 171968 460294 172020 460300
rect 171876 459944 171928 459950
rect 171876 459886 171928 459892
rect 171888 248334 171916 459886
rect 171980 248402 172008 460294
rect 172072 249286 172100 460362
rect 174450 459912 174506 459921
rect 174450 459847 174506 459856
rect 172152 456884 172204 456890
rect 172152 456826 172204 456832
rect 172060 249280 172112 249286
rect 172060 249222 172112 249228
rect 172164 249150 172192 456826
rect 172244 456340 172296 456346
rect 172244 456282 172296 456288
rect 172256 249218 172284 456282
rect 172336 454640 172388 454646
rect 172336 454582 172388 454588
rect 172348 349450 172376 454582
rect 172336 349444 172388 349450
rect 172336 349386 172388 349392
rect 174464 249762 174492 459847
rect 174452 249756 174504 249762
rect 174452 249698 174504 249704
rect 172244 249212 172296 249218
rect 172244 249154 172296 249160
rect 172152 249144 172204 249150
rect 172152 249086 172204 249092
rect 171968 248396 172020 248402
rect 171968 248338 172020 248344
rect 171876 248328 171928 248334
rect 171876 248270 171928 248276
rect 174556 248033 174584 462538
rect 174648 248878 174676 463286
rect 177304 461984 177356 461990
rect 177304 461926 177356 461932
rect 174820 461440 174872 461446
rect 174820 461382 174872 461388
rect 174728 461304 174780 461310
rect 174728 461246 174780 461252
rect 174740 249014 174768 461246
rect 174832 249558 174860 461382
rect 174912 461372 174964 461378
rect 174912 461314 174964 461320
rect 174924 249694 174952 461314
rect 175186 460048 175242 460057
rect 175186 459983 175242 459992
rect 175002 459776 175058 459785
rect 175002 459711 175058 459720
rect 174912 249688 174964 249694
rect 174912 249630 174964 249636
rect 174820 249552 174872 249558
rect 174820 249494 174872 249500
rect 174728 249008 174780 249014
rect 174728 248950 174780 248956
rect 175016 248946 175044 459711
rect 175096 453688 175148 453694
rect 175096 453630 175148 453636
rect 175108 349081 175136 453630
rect 175094 349072 175150 349081
rect 175094 349007 175150 349016
rect 175200 249626 175228 459983
rect 177212 453212 177264 453218
rect 177212 453154 177264 453160
rect 177224 348362 177252 453154
rect 177212 348356 177264 348362
rect 177212 348298 177264 348304
rect 175188 249620 175240 249626
rect 175188 249562 175240 249568
rect 175004 248940 175056 248946
rect 175004 248882 175056 248888
rect 174636 248872 174688 248878
rect 174636 248814 174688 248820
rect 174542 248024 174598 248033
rect 174542 247959 174598 247968
rect 171782 247888 171838 247897
rect 171782 247823 171838 247832
rect 177316 247722 177344 461926
rect 195980 461848 196032 461854
rect 195980 461790 196032 461796
rect 177488 461508 177540 461514
rect 177488 461450 177540 461456
rect 177396 460624 177448 460630
rect 177396 460566 177448 460572
rect 177304 247716 177356 247722
rect 177304 247658 177356 247664
rect 177408 247518 177436 460566
rect 177500 249422 177528 461450
rect 183006 461408 183062 461417
rect 183006 461343 183062 461352
rect 182822 461272 182878 461281
rect 182822 461207 182878 461216
rect 177672 460080 177724 460086
rect 177672 460022 177724 460028
rect 177580 458380 177632 458386
rect 177580 458322 177632 458328
rect 177488 249416 177540 249422
rect 177488 249358 177540 249364
rect 177592 247790 177620 458322
rect 177684 249354 177712 460022
rect 180616 457904 180668 457910
rect 180616 457846 180668 457852
rect 180062 457736 180118 457745
rect 180062 457671 180118 457680
rect 180432 457700 180484 457706
rect 179972 453280 180024 453286
rect 179972 453222 180024 453228
rect 177948 450764 178000 450770
rect 177948 450706 178000 450712
rect 177856 450220 177908 450226
rect 177856 450162 177908 450168
rect 177762 448760 177818 448769
rect 177762 448695 177818 448704
rect 177672 249348 177724 249354
rect 177672 249290 177724 249296
rect 177776 247858 177804 448695
rect 177868 249490 177896 450162
rect 177856 249484 177908 249490
rect 177856 249426 177908 249432
rect 177960 249082 177988 450706
rect 179984 347206 180012 453222
rect 179972 347200 180024 347206
rect 179972 347142 180024 347148
rect 177948 249076 178000 249082
rect 177948 249018 178000 249024
rect 177764 247852 177816 247858
rect 177764 247794 177816 247800
rect 177580 247784 177632 247790
rect 177580 247726 177632 247732
rect 177396 247512 177448 247518
rect 177396 247454 177448 247460
rect 179420 240780 179472 240786
rect 179420 240722 179472 240728
rect 172520 228404 172572 228410
rect 172520 228346 172572 228352
rect 170496 20664 170548 20670
rect 170496 20606 170548 20612
rect 172532 16574 172560 228346
rect 176660 227044 176712 227050
rect 176660 226986 176712 226992
rect 172532 16546 172744 16574
rect 170404 6860 170456 6866
rect 170404 6802 170456 6808
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 176672 480 176700 226986
rect 179432 16574 179460 240722
rect 180076 147558 180104 457671
rect 180432 457642 180484 457648
rect 180340 457564 180392 457570
rect 180340 457506 180392 457512
rect 180248 457428 180300 457434
rect 180248 457370 180300 457376
rect 180156 457360 180208 457366
rect 180156 457302 180208 457308
rect 180064 147552 180116 147558
rect 180064 147494 180116 147500
rect 180168 147393 180196 457302
rect 180260 148646 180288 457370
rect 180248 148640 180300 148646
rect 180248 148582 180300 148588
rect 180352 148578 180380 457506
rect 180444 247926 180472 457642
rect 180524 457020 180576 457026
rect 180524 456962 180576 456968
rect 180536 248266 180564 456962
rect 180524 248260 180576 248266
rect 180524 248202 180576 248208
rect 180628 248130 180656 457846
rect 182732 453348 182784 453354
rect 182732 453290 182784 453296
rect 180706 451752 180762 451761
rect 180706 451687 180762 451696
rect 180720 248169 180748 451687
rect 182744 348838 182772 453290
rect 182732 348832 182784 348838
rect 182732 348774 182784 348780
rect 180706 248160 180762 248169
rect 180616 248124 180668 248130
rect 180706 248095 180762 248104
rect 180616 248066 180668 248072
rect 180432 247920 180484 247926
rect 180432 247862 180484 247868
rect 180340 148572 180392 148578
rect 180340 148514 180392 148520
rect 182836 148170 182864 461207
rect 182914 457192 182970 457201
rect 182914 457127 182970 457136
rect 182824 148164 182876 148170
rect 182824 148106 182876 148112
rect 180154 147384 180210 147393
rect 180154 147319 180210 147328
rect 182928 146946 182956 457127
rect 183020 148238 183048 461343
rect 183190 461136 183246 461145
rect 183190 461071 183246 461080
rect 183098 459232 183154 459241
rect 183098 459167 183154 459176
rect 183112 148306 183140 459167
rect 183204 149025 183232 461071
rect 183374 461000 183430 461009
rect 183374 460935 183430 460944
rect 183284 457632 183336 457638
rect 183284 457574 183336 457580
rect 183190 149016 183246 149025
rect 183190 148951 183246 148960
rect 183296 148510 183324 457574
rect 183388 148889 183416 460935
rect 185676 459332 185728 459338
rect 185676 459274 185728 459280
rect 185582 458688 185638 458697
rect 185582 458623 185638 458632
rect 183466 450256 183522 450265
rect 183466 450191 183522 450200
rect 183480 149054 183508 450191
rect 184204 434036 184256 434042
rect 184204 433978 184256 433984
rect 184216 248402 184244 433978
rect 184204 248396 184256 248402
rect 184204 248338 184256 248344
rect 183560 225616 183612 225622
rect 183560 225558 183612 225564
rect 183468 149048 183520 149054
rect 183468 148990 183520 148996
rect 183374 148880 183430 148889
rect 183374 148815 183430 148824
rect 183284 148504 183336 148510
rect 183284 148446 183336 148452
rect 183100 148300 183152 148306
rect 183100 148242 183152 148248
rect 183008 148232 183060 148238
rect 183008 148174 183060 148180
rect 182916 146940 182968 146946
rect 182916 146882 182968 146888
rect 183572 16574 183600 225558
rect 185596 147286 185624 458623
rect 185688 148918 185716 459274
rect 188528 459264 188580 459270
rect 188528 459206 188580 459212
rect 185766 459096 185822 459105
rect 185766 459031 185822 459040
rect 185676 148912 185728 148918
rect 185676 148854 185728 148860
rect 185584 147280 185636 147286
rect 185584 147222 185636 147228
rect 185780 147082 185808 459031
rect 185950 458552 186006 458561
rect 185950 458487 186006 458496
rect 188344 458516 188396 458522
rect 185858 454064 185914 454073
rect 185858 453999 185914 454008
rect 185872 148442 185900 453999
rect 185964 148986 185992 458487
rect 188344 458458 188396 458464
rect 186964 458448 187016 458454
rect 186964 458390 187016 458396
rect 186136 450492 186188 450498
rect 186136 450434 186188 450440
rect 186044 450356 186096 450362
rect 186044 450298 186096 450304
rect 185952 148980 186004 148986
rect 185952 148922 186004 148928
rect 185860 148436 185912 148442
rect 185860 148378 185912 148384
rect 186056 147354 186084 450298
rect 186148 347342 186176 450434
rect 186976 347750 187004 458390
rect 187056 458312 187108 458318
rect 187056 458254 187108 458260
rect 186964 347744 187016 347750
rect 186964 347686 187016 347692
rect 187068 347614 187096 458254
rect 187514 452160 187570 452169
rect 187514 452095 187570 452104
rect 188252 452124 188304 452130
rect 187422 449576 187478 449585
rect 187422 449511 187478 449520
rect 187056 347608 187108 347614
rect 187056 347550 187108 347556
rect 186136 347336 186188 347342
rect 186136 347278 186188 347284
rect 186320 242208 186372 242214
rect 186320 242150 186372 242156
rect 186044 147348 186096 147354
rect 186044 147290 186096 147296
rect 185768 147076 185820 147082
rect 185768 147018 185820 147024
rect 186332 16574 186360 242150
rect 187436 134570 187464 449511
rect 187528 134706 187556 452095
rect 188252 452066 188304 452072
rect 187608 451308 187660 451314
rect 187608 451250 187660 451256
rect 187516 134700 187568 134706
rect 187516 134642 187568 134648
rect 187620 134638 187648 451250
rect 188264 349178 188292 452066
rect 188252 349172 188304 349178
rect 188252 349114 188304 349120
rect 188356 147422 188384 458458
rect 188434 457056 188490 457065
rect 188434 456991 188490 457000
rect 188448 147490 188476 456991
rect 188540 148714 188568 459206
rect 188896 458924 188948 458930
rect 188896 458866 188948 458872
rect 188620 458584 188672 458590
rect 188620 458526 188672 458532
rect 188632 148782 188660 458526
rect 188710 456920 188766 456929
rect 188710 456855 188766 456864
rect 188724 148850 188752 456855
rect 188804 456204 188856 456210
rect 188804 456146 188856 456152
rect 188712 148844 188764 148850
rect 188712 148786 188764 148792
rect 188620 148776 188672 148782
rect 188620 148718 188672 148724
rect 188528 148708 188580 148714
rect 188528 148650 188580 148656
rect 188816 148374 188844 456146
rect 188908 347682 188936 458866
rect 191196 455864 191248 455870
rect 191196 455806 191248 455812
rect 188988 454980 189040 454986
rect 188988 454922 189040 454928
rect 188896 347676 188948 347682
rect 188896 347618 188948 347624
rect 189000 346390 189028 454922
rect 189816 453416 189868 453422
rect 189816 453358 189868 453364
rect 189722 453248 189778 453257
rect 189722 453183 189778 453192
rect 188988 346384 189040 346390
rect 188988 346326 189040 346332
rect 188804 148368 188856 148374
rect 188804 148310 188856 148316
rect 189736 147626 189764 453183
rect 189828 347410 189856 453358
rect 190274 452432 190330 452441
rect 190274 452367 190330 452376
rect 189908 451988 189960 451994
rect 189908 451930 189960 451936
rect 189920 348498 189948 451930
rect 190000 451920 190052 451926
rect 190000 451862 190052 451868
rect 190012 349246 190040 451862
rect 190182 450664 190238 450673
rect 190182 450599 190238 450608
rect 190000 349240 190052 349246
rect 190000 349182 190052 349188
rect 189908 348492 189960 348498
rect 189908 348434 189960 348440
rect 189816 347404 189868 347410
rect 189816 347346 189868 347352
rect 190196 238066 190224 450599
rect 190184 238060 190236 238066
rect 190184 238002 190236 238008
rect 189724 147620 189776 147626
rect 189724 147562 189776 147568
rect 188436 147484 188488 147490
rect 188436 147426 188488 147432
rect 188344 147416 188396 147422
rect 188344 147358 188396 147364
rect 187608 134632 187660 134638
rect 187608 134574 187660 134580
rect 187424 134564 187476 134570
rect 187424 134506 187476 134512
rect 190288 46918 190316 452367
rect 191012 452056 191064 452062
rect 191012 451998 191064 452004
rect 190920 451648 190972 451654
rect 190920 451590 190972 451596
rect 190366 451480 190422 451489
rect 190366 451415 190422 451424
rect 190276 46912 190328 46918
rect 190276 46854 190328 46860
rect 179432 16546 180288 16574
rect 183572 16546 183784 16574
rect 186332 16546 186912 16574
rect 180260 480 180288 16546
rect 183756 480 183784 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 190380 6866 190408 451415
rect 190828 449880 190880 449886
rect 190828 449822 190880 449828
rect 190840 449546 190868 449822
rect 190828 449540 190880 449546
rect 190828 449482 190880 449488
rect 190932 349314 190960 451590
rect 190920 349308 190972 349314
rect 190920 349250 190972 349256
rect 190826 348664 190882 348673
rect 190826 348599 190882 348608
rect 190840 348566 190868 348599
rect 190828 348560 190880 348566
rect 191024 348514 191052 451998
rect 191102 450936 191158 450945
rect 191102 450871 191158 450880
rect 190828 348502 190880 348508
rect 190932 348486 191052 348514
rect 190932 348430 190960 348486
rect 190920 348424 190972 348430
rect 190920 348366 190972 348372
rect 191116 347698 191144 450871
rect 190748 347670 191144 347698
rect 190642 347440 190698 347449
rect 190642 347375 190698 347384
rect 190656 347177 190684 347375
rect 190642 347168 190698 347177
rect 190642 347103 190698 347112
rect 190748 345014 190776 347670
rect 190826 347576 190882 347585
rect 191208 347562 191236 455806
rect 191288 454844 191340 454850
rect 191288 454786 191340 454792
rect 191300 347585 191328 454786
rect 195992 454034 196020 461790
rect 196084 458844 196112 466482
rect 196164 466472 196216 466478
rect 196164 466414 196216 466420
rect 196176 461854 196204 466414
rect 197452 465180 197504 465186
rect 197452 465122 197504 465128
rect 196164 461848 196216 461854
rect 196164 461790 196216 461796
rect 197360 458856 197412 458862
rect 196084 458816 196296 458844
rect 196268 454034 196296 458816
rect 197360 458798 197412 458804
rect 195992 454006 196204 454034
rect 196268 454006 196388 454034
rect 191472 453484 191524 453490
rect 191472 453426 191524 453432
rect 191380 453144 191432 453150
rect 191380 453086 191432 453092
rect 190826 347511 190828 347520
rect 190880 347511 190882 347520
rect 190932 347534 191236 347562
rect 191286 347576 191342 347585
rect 190828 347482 190880 347488
rect 190932 347478 190960 347534
rect 191286 347511 191342 347520
rect 190920 347472 190972 347478
rect 190826 347440 190882 347449
rect 190920 347414 190972 347420
rect 190826 347375 190882 347384
rect 190840 347274 190868 347375
rect 190828 347268 190880 347274
rect 190828 347210 190880 347216
rect 191392 347154 191420 453086
rect 191484 347313 191512 453426
rect 195150 452704 195206 452713
rect 193864 452668 193916 452674
rect 195150 452639 195206 452648
rect 193864 452610 193916 452616
rect 193218 451888 193274 451897
rect 191748 451852 191800 451858
rect 193218 451823 193274 451832
rect 191748 451794 191800 451800
rect 191656 450832 191708 450838
rect 191656 450774 191708 450780
rect 191564 450424 191616 450430
rect 191564 450366 191616 450372
rect 191576 347449 191604 450366
rect 191668 347721 191696 450774
rect 191760 348673 191788 451794
rect 191840 450288 191892 450294
rect 191840 450230 191892 450236
rect 191746 348664 191802 348673
rect 191746 348599 191802 348608
rect 191654 347712 191710 347721
rect 191654 347647 191710 347656
rect 191562 347440 191618 347449
rect 191562 347375 191618 347384
rect 191470 347304 191526 347313
rect 191470 347239 191526 347248
rect 190932 347138 191420 347154
rect 190920 347132 191420 347138
rect 190972 347126 191420 347132
rect 190920 347074 190972 347080
rect 191852 345137 191880 450230
rect 193232 449834 193260 451823
rect 193678 451480 193734 451489
rect 193678 451415 193734 451424
rect 193692 449956 193720 451415
rect 193876 449886 193904 452610
rect 194782 452432 194838 452441
rect 194782 452367 194838 452376
rect 194138 450392 194194 450401
rect 194138 450327 194194 450336
rect 194152 449970 194180 450327
rect 194152 449942 194442 449970
rect 194796 449956 194824 452367
rect 195164 449956 195192 452639
rect 195886 452160 195942 452169
rect 195886 452095 195942 452104
rect 195900 449956 195928 452095
rect 196176 449970 196204 454006
rect 196360 449970 196388 454006
rect 196992 451308 197044 451314
rect 196992 451250 197044 451256
rect 196176 449942 196282 449970
rect 196360 449942 196650 449970
rect 197004 449956 197032 451250
rect 197372 449956 197400 458798
rect 197464 456906 197492 465122
rect 197544 465112 197596 465118
rect 197544 465054 197596 465060
rect 197556 458862 197584 465054
rect 197544 458856 197596 458862
rect 197544 458798 197596 458804
rect 197464 456878 197584 456906
rect 197556 454034 197584 456878
rect 197648 456794 197676 466550
rect 198016 458998 198044 682382
rect 198096 682372 198148 682378
rect 198096 682314 198148 682320
rect 198108 459066 198136 682314
rect 198200 459134 198228 682518
rect 198280 682508 198332 682514
rect 198280 682450 198332 682456
rect 198188 459128 198240 459134
rect 198188 459070 198240 459076
rect 198096 459060 198148 459066
rect 198096 459002 198148 459008
rect 198004 458992 198056 458998
rect 198004 458934 198056 458940
rect 198292 458862 198320 682450
rect 198372 681760 198424 681766
rect 198372 681702 198424 681708
rect 198384 460290 198412 681702
rect 198924 466880 198976 466886
rect 198924 466822 198976 466828
rect 198832 466812 198884 466818
rect 198832 466754 198884 466760
rect 198740 466744 198792 466750
rect 198740 466686 198792 466692
rect 198372 460284 198424 460290
rect 198372 460226 198424 460232
rect 198280 458856 198332 458862
rect 198280 458798 198332 458804
rect 197648 456766 198228 456794
rect 197464 454006 197584 454034
rect 197464 449970 197492 454006
rect 197818 450664 197874 450673
rect 197818 450599 197874 450608
rect 197832 449970 197860 450599
rect 198200 449970 198228 456766
rect 198752 452742 198780 466686
rect 198740 452736 198792 452742
rect 198740 452678 198792 452684
rect 198844 452606 198872 466754
rect 198832 452600 198884 452606
rect 198832 452542 198884 452548
rect 198936 449970 198964 466822
rect 199396 464506 199424 700334
rect 202144 683188 202196 683194
rect 202144 683130 202196 683136
rect 200120 466676 200172 466682
rect 200120 466618 200172 466624
rect 199384 464500 199436 464506
rect 199384 464442 199436 464448
rect 199016 463752 199068 463758
rect 199016 463694 199068 463700
rect 197464 449942 197754 449970
rect 197832 449942 198122 449970
rect 198200 449942 198490 449970
rect 198858 449942 198964 449970
rect 199028 449970 199056 463694
rect 199292 452736 199344 452742
rect 199292 452678 199344 452684
rect 199304 449970 199332 452678
rect 199660 452600 199712 452606
rect 199660 452542 199712 452548
rect 199672 449970 199700 452542
rect 200132 449970 200160 466618
rect 202156 463282 202184 683130
rect 202144 463276 202196 463282
rect 202144 463218 202196 463224
rect 203536 461854 203564 700334
rect 206284 700324 206336 700330
rect 206284 700266 206336 700272
rect 212540 700324 212592 700330
rect 212540 700266 212592 700272
rect 205640 498840 205692 498846
rect 205640 498782 205692 498788
rect 204260 470620 204312 470626
rect 204260 470562 204312 470568
rect 203524 461848 203576 461854
rect 203524 461790 203576 461796
rect 202880 461168 202932 461174
rect 202880 461110 202932 461116
rect 201500 461100 201552 461106
rect 201500 461042 201552 461048
rect 200764 456136 200816 456142
rect 200764 456078 200816 456084
rect 200776 455870 200804 456078
rect 200764 455864 200816 455870
rect 200764 455806 200816 455812
rect 200670 454880 200726 454889
rect 200670 454815 200726 454824
rect 199028 449942 199226 449970
rect 199304 449942 199594 449970
rect 199672 449942 199962 449970
rect 200132 449942 200330 449970
rect 200684 449956 200712 454815
rect 201406 454336 201462 454345
rect 201406 454271 201462 454280
rect 201038 454200 201094 454209
rect 201038 454135 201094 454144
rect 201052 449956 201080 454135
rect 201420 449956 201448 454271
rect 201512 449970 201540 461042
rect 202510 456240 202566 456249
rect 202510 456175 202566 456184
rect 202142 454472 202198 454481
rect 202142 454407 202198 454416
rect 201512 449942 201802 449970
rect 202156 449956 202184 454407
rect 202524 449956 202552 456175
rect 202892 452742 202920 461110
rect 202972 461032 203024 461038
rect 202972 460974 203024 460980
rect 202880 452736 202932 452742
rect 202880 452678 202932 452684
rect 202984 449970 203012 460974
rect 203064 460964 203116 460970
rect 203064 460906 203116 460912
rect 202906 449942 203012 449970
rect 203076 449970 203104 460906
rect 203338 459640 203394 459649
rect 203338 459575 203394 459584
rect 203352 449970 203380 459575
rect 203708 452736 203760 452742
rect 203708 452678 203760 452684
rect 203720 449970 203748 452678
rect 204272 452606 204300 470562
rect 204352 468580 204404 468586
rect 204352 468522 204404 468528
rect 204364 452742 204392 468522
rect 204444 461236 204496 461242
rect 204444 461178 204496 461184
rect 204352 452736 204404 452742
rect 204352 452678 204404 452684
rect 204260 452600 204312 452606
rect 204260 452542 204312 452548
rect 204456 449970 204484 461178
rect 204536 459604 204588 459610
rect 204536 459546 204588 459552
rect 203076 449942 203274 449970
rect 203352 449942 203642 449970
rect 203720 449942 204010 449970
rect 204378 449942 204484 449970
rect 204548 449970 204576 459546
rect 204812 452736 204864 452742
rect 204812 452678 204864 452684
rect 204824 449970 204852 452678
rect 205180 452600 205232 452606
rect 205180 452542 205232 452548
rect 205192 449970 205220 452542
rect 205652 449970 205680 498782
rect 205732 489184 205784 489190
rect 205732 489126 205784 489132
rect 205744 452606 205772 489126
rect 205824 479528 205876 479534
rect 205824 479470 205876 479476
rect 205836 452742 205864 479470
rect 206296 476950 206324 700266
rect 208400 630692 208452 630698
rect 208400 630634 208452 630640
rect 207020 480956 207072 480962
rect 207020 480898 207072 480904
rect 206284 476944 206336 476950
rect 206284 476886 206336 476892
rect 205916 474020 205968 474026
rect 205916 473962 205968 473968
rect 205824 452736 205876 452742
rect 205824 452678 205876 452684
rect 205732 452600 205784 452606
rect 205732 452542 205784 452548
rect 205928 449970 205956 473962
rect 207032 452742 207060 480898
rect 207112 469940 207164 469946
rect 207112 469882 207164 469888
rect 207124 456794 207152 469882
rect 207204 461712 207256 461718
rect 207204 461654 207256 461660
rect 207216 460934 207244 461654
rect 207216 460906 207796 460934
rect 207124 456766 207244 456794
rect 206284 452736 206336 452742
rect 206284 452678 206336 452684
rect 207020 452736 207072 452742
rect 207020 452678 207072 452684
rect 206296 449970 206324 452678
rect 206652 452600 206704 452606
rect 206652 452542 206704 452548
rect 206664 449970 206692 452542
rect 207216 449970 207244 456766
rect 207388 452736 207440 452742
rect 207388 452678 207440 452684
rect 207400 449970 207428 452678
rect 207768 449970 207796 460906
rect 208308 451580 208360 451586
rect 208308 451522 208360 451528
rect 208320 449970 208348 451522
rect 208412 450378 208440 630634
rect 209780 588600 209832 588606
rect 209780 588542 209832 588548
rect 208492 478236 208544 478242
rect 208492 478178 208544 478184
rect 208504 452742 208532 478178
rect 208584 467220 208636 467226
rect 208584 467162 208636 467168
rect 208492 452736 208544 452742
rect 208492 452678 208544 452684
rect 208596 451586 208624 467162
rect 208676 464432 208728 464438
rect 208676 464374 208728 464380
rect 208688 460934 208716 464374
rect 208688 460906 208900 460934
rect 208584 451580 208636 451586
rect 208584 451522 208636 451528
rect 208412 450350 208532 450378
rect 208504 449970 208532 450350
rect 208872 449970 208900 460906
rect 209228 452736 209280 452742
rect 209228 452678 209280 452684
rect 209240 449970 209268 452678
rect 209792 452606 209820 588542
rect 211160 587172 211212 587178
rect 211160 587114 211212 587120
rect 209872 585812 209924 585818
rect 209872 585754 209924 585760
rect 209884 452742 209912 585754
rect 209964 482384 210016 482390
rect 209964 482326 210016 482332
rect 209872 452736 209924 452742
rect 209872 452678 209924 452684
rect 209780 452600 209832 452606
rect 209780 452542 209832 452548
rect 209976 449970 210004 482326
rect 210056 465724 210108 465730
rect 210056 465666 210108 465672
rect 204548 449942 204746 449970
rect 204824 449942 205114 449970
rect 205192 449942 205482 449970
rect 205652 449942 205850 449970
rect 205928 449942 206218 449970
rect 206296 449942 206586 449970
rect 206664 449942 206954 449970
rect 207216 449942 207322 449970
rect 207400 449942 207690 449970
rect 207768 449942 208058 449970
rect 208320 449942 208426 449970
rect 208504 449942 208794 449970
rect 208872 449942 209162 449970
rect 209240 449942 209530 449970
rect 209898 449942 210004 449970
rect 210068 449970 210096 465666
rect 211172 452742 211200 587114
rect 211252 584452 211304 584458
rect 211252 584394 211304 584400
rect 210332 452736 210384 452742
rect 210332 452678 210384 452684
rect 211160 452736 211212 452742
rect 211160 452678 211212 452684
rect 210344 449970 210372 452678
rect 210700 452600 210752 452606
rect 210700 452542 210752 452548
rect 210516 451308 210568 451314
rect 210516 451250 210568 451256
rect 210424 450900 210476 450906
rect 210424 450842 210476 450848
rect 210436 450537 210464 450842
rect 210528 450634 210556 451250
rect 210516 450628 210568 450634
rect 210516 450570 210568 450576
rect 210422 450528 210478 450537
rect 210422 450463 210478 450472
rect 210712 449970 210740 452542
rect 211264 449970 211292 584394
rect 211344 505776 211396 505782
rect 211344 505718 211396 505724
rect 211356 456794 211384 505718
rect 211436 500268 211488 500274
rect 211436 500210 211488 500216
rect 211448 460934 211476 500210
rect 211448 460906 212212 460934
rect 211356 456766 211844 456794
rect 211436 452736 211488 452742
rect 211436 452678 211488 452684
rect 211448 449970 211476 452678
rect 211816 449970 211844 456766
rect 212184 449970 212212 460906
rect 212552 452742 212580 700266
rect 218992 697610 219020 703520
rect 215300 697604 215352 697610
rect 215300 697546 215352 697552
rect 218980 697604 219032 697610
rect 218980 697546 219032 697552
rect 213920 507136 213972 507142
rect 213920 507078 213972 507084
rect 212632 502988 212684 502994
rect 212632 502930 212684 502936
rect 212540 452736 212592 452742
rect 212540 452678 212592 452684
rect 212644 452606 212672 502930
rect 212724 501628 212776 501634
rect 212724 501570 212776 501576
rect 212632 452600 212684 452606
rect 212632 452542 212684 452548
rect 212736 449970 212764 501570
rect 213932 452742 213960 507078
rect 214012 504416 214064 504422
rect 214012 504358 214064 504364
rect 212908 452736 212960 452742
rect 212908 452678 212960 452684
rect 213920 452736 213972 452742
rect 213920 452678 213972 452684
rect 212920 449970 212948 452678
rect 213276 452600 213328 452606
rect 213276 452542 213328 452548
rect 213288 449970 213316 452542
rect 214024 449970 214052 504358
rect 214104 476876 214156 476882
rect 214104 476818 214156 476824
rect 214116 453558 214144 476818
rect 214196 472728 214248 472734
rect 214196 472670 214248 472676
rect 214208 460934 214236 472670
rect 214208 460906 214420 460934
rect 214104 453552 214156 453558
rect 214104 453494 214156 453500
rect 214104 452736 214156 452742
rect 214104 452678 214156 452684
rect 210068 449942 210266 449970
rect 210344 449942 210634 449970
rect 210712 449942 211002 449970
rect 211264 449942 211370 449970
rect 211448 449942 211738 449970
rect 211816 449942 212106 449970
rect 212184 449942 212474 449970
rect 212736 449942 212842 449970
rect 212920 449942 213210 449970
rect 213288 449942 213578 449970
rect 213946 449942 214052 449970
rect 214116 449970 214144 452678
rect 214392 449970 214420 460906
rect 215312 456006 215340 697546
rect 219440 692096 219492 692102
rect 219440 692038 219492 692044
rect 218060 690668 218112 690674
rect 218060 690610 218112 690616
rect 216680 689308 216732 689314
rect 216680 689250 216732 689256
rect 215392 492040 215444 492046
rect 215392 491982 215444 491988
rect 215300 456000 215352 456006
rect 215300 455942 215352 455948
rect 214748 453552 214800 453558
rect 214748 453494 214800 453500
rect 214760 449970 214788 453494
rect 214116 449942 214314 449970
rect 214392 449942 214682 449970
rect 214760 449942 215050 449970
rect 215404 449956 215432 491982
rect 215576 461848 215628 461854
rect 215576 461790 215628 461796
rect 215484 461644 215536 461650
rect 215484 461586 215536 461592
rect 215496 449970 215524 461586
rect 215588 460934 215616 461790
rect 215588 460906 215892 460934
rect 215864 449970 215892 460906
rect 216692 456550 216720 689250
rect 216772 686520 216824 686526
rect 216772 686462 216824 686468
rect 216784 458658 216812 686462
rect 216864 685160 216916 685166
rect 216864 685102 216916 685108
rect 216772 458652 216824 458658
rect 216772 458594 216824 458600
rect 216680 456544 216732 456550
rect 216680 456486 216732 456492
rect 216876 456226 216904 685102
rect 216956 464500 217008 464506
rect 216956 464442 217008 464448
rect 216968 460934 216996 464442
rect 216968 460906 217364 460934
rect 216956 456544 217008 456550
rect 216956 456486 217008 456492
rect 216692 456198 216904 456226
rect 216220 456000 216272 456006
rect 216220 455942 216272 455948
rect 216232 449970 216260 455942
rect 216692 449970 216720 456198
rect 216968 455954 216996 456486
rect 216784 455926 216996 455954
rect 216784 450242 216812 455926
rect 216784 450214 216996 450242
rect 216968 449970 216996 450214
rect 217336 449970 217364 460906
rect 217692 458652 217744 458658
rect 217692 458594 217744 458600
rect 217704 449970 217732 458594
rect 218072 449970 218100 690610
rect 218152 687948 218204 687954
rect 218152 687890 218204 687896
rect 218164 456006 218192 687890
rect 218244 476944 218296 476950
rect 218244 476886 218296 476892
rect 218256 460934 218284 476886
rect 218256 460906 218468 460934
rect 218152 456000 218204 456006
rect 218152 455942 218204 455948
rect 218440 449970 218468 460906
rect 219452 456550 219480 692038
rect 224224 683188 224276 683194
rect 224224 683130 224276 683136
rect 222844 616888 222896 616894
rect 222844 616830 222896 616836
rect 222200 481024 222252 481030
rect 222200 480966 222252 480972
rect 220820 479596 220872 479602
rect 220820 479538 220872 479544
rect 219532 469872 219584 469878
rect 219532 469814 219584 469820
rect 219544 458658 219572 469814
rect 219624 468512 219676 468518
rect 219624 468454 219676 468460
rect 219532 458652 219584 458658
rect 219532 458594 219584 458600
rect 219440 456544 219492 456550
rect 219440 456486 219492 456492
rect 219636 456090 219664 468454
rect 219716 463276 219768 463282
rect 219716 463218 219768 463224
rect 219728 460934 219756 463218
rect 219728 460906 219940 460934
rect 219716 456544 219768 456550
rect 219716 456486 219768 456492
rect 219452 456062 219664 456090
rect 218796 456000 218848 456006
rect 218796 455942 218848 455948
rect 218808 449970 218836 455942
rect 215496 449942 215786 449970
rect 215864 449942 216154 449970
rect 216232 449942 216522 449970
rect 216692 449942 216890 449970
rect 216968 449942 217258 449970
rect 217336 449942 217626 449970
rect 217704 449942 217994 449970
rect 218072 449942 218362 449970
rect 218440 449942 218730 449970
rect 218808 449942 219098 449970
rect 219452 449956 219480 456062
rect 219728 455818 219756 456486
rect 219544 455790 219756 455818
rect 219544 449970 219572 455790
rect 219912 449970 219940 460906
rect 220268 458652 220320 458658
rect 220268 458594 220320 458600
rect 220280 449970 220308 458594
rect 220832 456006 220860 479538
rect 220912 478168 220964 478174
rect 220912 478110 220964 478116
rect 220820 456000 220872 456006
rect 220820 455942 220872 455948
rect 219544 449942 219834 449970
rect 219912 449942 220202 449970
rect 220280 449942 220570 449970
rect 220924 449956 220952 478110
rect 221004 471300 221056 471306
rect 221004 471242 221056 471248
rect 221016 458726 221044 471242
rect 221096 464364 221148 464370
rect 221096 464306 221148 464312
rect 221004 458720 221056 458726
rect 221004 458662 221056 458668
rect 221108 449970 221136 464306
rect 221372 458720 221424 458726
rect 221372 458662 221424 458668
rect 221384 449970 221412 458662
rect 221740 456000 221792 456006
rect 221740 455942 221792 455948
rect 221752 449970 221780 455942
rect 222212 450294 222240 480966
rect 222292 472660 222344 472666
rect 222292 472602 222344 472608
rect 222304 455682 222332 472602
rect 222384 467152 222436 467158
rect 222384 467094 222436 467100
rect 222396 456006 222424 467094
rect 222476 465792 222528 465798
rect 222476 465734 222528 465740
rect 222488 460934 222516 465734
rect 222856 461718 222884 616830
rect 224236 482390 224264 683130
rect 231124 670744 231176 670750
rect 231124 670686 231176 670692
rect 228364 590708 228416 590714
rect 228364 590650 228416 590656
rect 226984 484424 227036 484430
rect 226984 484366 227036 484372
rect 224224 482384 224276 482390
rect 224224 482326 224276 482332
rect 223580 482316 223632 482322
rect 223580 482258 223632 482264
rect 222844 461712 222896 461718
rect 222844 461654 222896 461660
rect 222488 460906 222700 460934
rect 222384 456000 222436 456006
rect 222384 455942 222436 455948
rect 222304 455654 222608 455682
rect 222476 451308 222528 451314
rect 222476 451250 222528 451256
rect 222108 450288 222160 450294
rect 222108 450230 222160 450236
rect 222200 450288 222252 450294
rect 222200 450230 222252 450236
rect 222120 450106 222148 450230
rect 222292 450152 222344 450158
rect 222120 450100 222292 450106
rect 222120 450094 222344 450100
rect 222120 450078 222332 450094
rect 222488 449970 222516 451250
rect 221108 449942 221306 449970
rect 221384 449942 221674 449970
rect 221752 449942 222042 449970
rect 222410 449942 222516 449970
rect 222580 449970 222608 455654
rect 222672 451314 222700 460906
rect 223212 456000 223264 456006
rect 223212 455942 223264 455948
rect 222660 451308 222712 451314
rect 222660 451250 222712 451256
rect 222844 450288 222896 450294
rect 222844 450230 222896 450236
rect 222856 449970 222884 450230
rect 223224 449970 223252 455942
rect 223592 450294 223620 482258
rect 223672 474768 223724 474774
rect 223672 474710 223724 474716
rect 223684 456006 223712 474710
rect 223764 474088 223816 474094
rect 223764 474030 223816 474036
rect 223672 456000 223724 456006
rect 223672 455942 223724 455948
rect 223580 450288 223632 450294
rect 223580 450230 223632 450236
rect 223776 449970 223804 474030
rect 226996 468586 227024 484366
rect 228376 469946 228404 590650
rect 228364 469940 228416 469946
rect 228364 469882 228416 469888
rect 226984 468580 227036 468586
rect 226984 468522 227036 468528
rect 231136 464438 231164 670686
rect 233884 643136 233936 643142
rect 233884 643078 233936 643084
rect 233896 467226 233924 643078
rect 233884 467220 233936 467226
rect 233884 467162 233936 467168
rect 231858 466576 231914 466585
rect 231858 466511 231914 466520
rect 231124 464432 231176 464438
rect 231124 464374 231176 464380
rect 225144 462392 225196 462398
rect 225144 462334 225196 462340
rect 224316 456000 224368 456006
rect 224316 455942 224368 455948
rect 223948 450288 224000 450294
rect 223948 450230 224000 450236
rect 223960 449970 223988 450230
rect 224328 449970 224356 455942
rect 224960 452668 225012 452674
rect 224960 452610 225012 452616
rect 222580 449942 222778 449970
rect 222856 449942 223146 449970
rect 223224 449942 223514 449970
rect 223776 449942 223882 449970
rect 223960 449942 224250 449970
rect 224328 449942 224618 449970
rect 224972 449956 225000 452610
rect 225156 449970 225184 462334
rect 229100 461916 229152 461922
rect 229100 461858 229152 461864
rect 226064 453008 226116 453014
rect 226064 452950 226116 452956
rect 225696 451308 225748 451314
rect 225696 451250 225748 451256
rect 225156 449942 225354 449970
rect 225708 449956 225736 451250
rect 226076 449956 226104 452950
rect 227536 452940 227588 452946
rect 227536 452882 227588 452888
rect 226432 452872 226484 452878
rect 226432 452814 226484 452820
rect 226444 449956 226472 452814
rect 227168 450152 227220 450158
rect 227168 450094 227220 450100
rect 226616 450016 226668 450022
rect 226668 449964 226826 449970
rect 226616 449958 226826 449964
rect 226628 449942 226826 449958
rect 227180 449956 227208 450094
rect 227548 449956 227576 452882
rect 229006 452840 229062 452849
rect 228640 452804 228692 452810
rect 229006 452775 229062 452784
rect 228640 452746 228692 452752
rect 227902 451888 227958 451897
rect 227902 451823 227958 451832
rect 227916 449956 227944 451823
rect 228652 449956 228680 452746
rect 229020 449956 229048 452775
rect 229112 449970 229140 461858
rect 231308 460488 231360 460494
rect 231308 460430 231360 460436
rect 230572 459876 230624 459882
rect 230572 459818 230624 459824
rect 230110 452024 230166 452033
rect 230110 451959 230166 451968
rect 229112 449942 229402 449970
rect 230124 449956 230152 451959
rect 230584 449970 230612 459818
rect 230664 458244 230716 458250
rect 230664 458186 230716 458192
rect 230506 449942 230612 449970
rect 230676 449970 230704 458186
rect 230940 454436 230992 454442
rect 230940 454378 230992 454384
rect 230952 449970 230980 454378
rect 231320 449970 231348 460430
rect 231872 449970 231900 466511
rect 231952 465248 232004 465254
rect 231952 465190 232004 465196
rect 231964 456006 231992 465190
rect 233516 463004 233568 463010
rect 233516 462946 233568 462952
rect 232044 462460 232096 462466
rect 232044 462402 232096 462408
rect 232056 460934 232084 462402
rect 232056 460906 232452 460934
rect 231952 456000 232004 456006
rect 231952 455942 232004 455948
rect 232318 449984 232374 449993
rect 230676 449942 230874 449970
rect 230952 449942 231242 449970
rect 231320 449942 231610 449970
rect 231872 449942 231978 449970
rect 232424 449970 232452 460906
rect 233332 459808 233384 459814
rect 233332 459750 233384 459756
rect 232780 456000 232832 456006
rect 232780 455942 232832 455948
rect 232792 449970 232820 455942
rect 233344 449970 233372 459750
rect 233528 449970 233556 462946
rect 234632 461650 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 249800 684956 249852 684962
rect 249800 684898 249852 684904
rect 248420 684888 248472 684894
rect 248420 684830 248472 684836
rect 244280 684820 244332 684826
rect 244280 684762 244332 684768
rect 242900 684752 242952 684758
rect 242900 684694 242952 684700
rect 240140 684684 240192 684690
rect 240140 684626 240192 684632
rect 238760 683596 238812 683602
rect 238760 683538 238812 683544
rect 237656 683528 237708 683534
rect 237656 683470 237708 683476
rect 236000 683460 236052 683466
rect 236000 683402 236052 683408
rect 234712 679448 234764 679454
rect 234712 679390 234764 679396
rect 234620 461644 234672 461650
rect 234620 461586 234672 461592
rect 234252 456272 234304 456278
rect 234252 456214 234304 456220
rect 233882 454744 233938 454753
rect 233882 454679 233938 454688
rect 233896 449970 233924 454679
rect 234264 449970 234292 456214
rect 234724 453014 234752 679390
rect 234802 461544 234858 461553
rect 234802 461479 234858 461488
rect 234712 453008 234764 453014
rect 234712 452950 234764 452956
rect 234816 449970 234844 461479
rect 234988 457496 235040 457502
rect 234988 457438 235040 457444
rect 235000 449970 235028 457438
rect 235356 453008 235408 453014
rect 235356 452950 235408 452956
rect 235368 449970 235396 452950
rect 232424 449942 232714 449970
rect 232792 449942 233082 449970
rect 233344 449942 233450 449970
rect 233528 449942 233818 449970
rect 233896 449942 234186 449970
rect 234264 449942 234554 449970
rect 234816 449942 234922 449970
rect 235000 449942 235290 449970
rect 235368 449942 235658 449970
rect 236012 449956 236040 683402
rect 236090 681048 236146 681057
rect 236090 680983 236146 680992
rect 236104 453014 236132 680983
rect 236184 680808 236236 680814
rect 236184 680750 236236 680756
rect 236092 453008 236144 453014
rect 236092 452950 236144 452956
rect 236196 452946 236224 680750
rect 237470 680368 237526 680377
rect 237470 680303 237526 680312
rect 236276 476808 236328 476814
rect 236276 476750 236328 476756
rect 236288 460934 236316 476750
rect 236288 460906 236500 460934
rect 236184 452940 236236 452946
rect 236184 452882 236236 452888
rect 236472 449970 236500 460906
rect 237380 459128 237432 459134
rect 237380 459070 237432 459076
rect 236552 453008 236604 453014
rect 236552 452950 236604 452956
rect 236394 449942 236500 449970
rect 236564 449970 236592 452950
rect 236828 452940 236880 452946
rect 236828 452882 236880 452888
rect 236840 449970 236868 452882
rect 237392 449970 237420 459070
rect 237484 453014 237512 680303
rect 237562 679552 237618 679561
rect 237562 679487 237618 679496
rect 237576 460834 237604 679487
rect 237564 460828 237616 460834
rect 237564 460770 237616 460776
rect 237472 453008 237524 453014
rect 237472 452950 237524 452956
rect 237668 449970 237696 683470
rect 237932 460828 237984 460834
rect 237932 460770 237984 460776
rect 237944 449970 237972 460770
rect 238300 453008 238352 453014
rect 238300 452950 238352 452956
rect 238312 449970 238340 452950
rect 238772 452946 238800 683538
rect 238852 683256 238904 683262
rect 238852 683198 238904 683204
rect 238760 452940 238812 452946
rect 238760 452882 238812 452888
rect 238864 452878 238892 683198
rect 238944 679380 238996 679386
rect 238944 679322 238996 679328
rect 238956 453014 238984 679322
rect 239036 679108 239088 679114
rect 239036 679050 239088 679056
rect 238944 453008 238996 453014
rect 238944 452950 238996 452956
rect 238852 452872 238904 452878
rect 238852 452814 238904 452820
rect 239048 449970 239076 679050
rect 240152 459542 240180 684626
rect 241520 684548 241572 684554
rect 241520 684490 241572 684496
rect 240230 680504 240286 680513
rect 240230 680439 240286 680448
rect 240140 459536 240192 459542
rect 240140 459478 240192 459484
rect 239128 453008 239180 453014
rect 239128 452950 239180 452956
rect 236564 449942 236762 449970
rect 236840 449942 237130 449970
rect 237392 449942 237498 449970
rect 237668 449942 237866 449970
rect 237944 449942 238234 449970
rect 238312 449942 238602 449970
rect 238970 449942 239076 449970
rect 239140 449970 239168 452950
rect 239404 452940 239456 452946
rect 239404 452882 239456 452888
rect 239416 449970 239444 452882
rect 239772 452872 239824 452878
rect 239772 452814 239824 452820
rect 239784 449970 239812 452814
rect 240244 449970 240272 680439
rect 240324 679176 240376 679182
rect 240324 679118 240376 679124
rect 240336 460934 240364 679118
rect 240336 460906 240548 460934
rect 240520 449970 240548 460906
rect 240876 459536 240928 459542
rect 240876 459478 240928 459484
rect 240888 449970 240916 459478
rect 241532 453014 241560 684490
rect 241612 683732 241664 683738
rect 241612 683674 241664 683680
rect 241520 453008 241572 453014
rect 241520 452950 241572 452956
rect 241624 449970 241652 683674
rect 241704 683324 241756 683330
rect 241704 683266 241756 683272
rect 239140 449942 239338 449970
rect 239416 449942 239706 449970
rect 239784 449942 240074 449970
rect 240244 449942 240442 449970
rect 240520 449942 240810 449970
rect 240888 449942 241178 449970
rect 241546 449942 241652 449970
rect 241716 449970 241744 683266
rect 241796 680400 241848 680406
rect 241796 680342 241848 680348
rect 241808 460934 241836 680342
rect 241808 460906 242020 460934
rect 241992 449970 242020 460906
rect 242348 453008 242400 453014
rect 242348 452950 242400 452956
rect 242360 449970 242388 452950
rect 242912 449970 242940 684694
rect 242992 684004 243044 684010
rect 242992 683946 243044 683952
rect 243004 453014 243032 683946
rect 243084 683800 243136 683806
rect 243084 683742 243136 683748
rect 242992 453008 243044 453014
rect 242992 452950 243044 452956
rect 243096 449970 243124 683742
rect 243176 681352 243228 681358
rect 243176 681294 243228 681300
rect 243188 460934 243216 681294
rect 243188 460906 243860 460934
rect 243452 453008 243504 453014
rect 243452 452950 243504 452956
rect 243464 449970 243492 452950
rect 243832 449970 243860 460906
rect 244292 456550 244320 684762
rect 245660 684072 245712 684078
rect 245660 684014 245712 684020
rect 244372 683664 244424 683670
rect 244372 683606 244424 683612
rect 244280 456544 244332 456550
rect 244280 456486 244332 456492
rect 244384 456006 244412 683606
rect 244462 682680 244518 682689
rect 244462 682615 244518 682624
rect 244372 456000 244424 456006
rect 244372 455942 244424 455948
rect 244476 450294 244504 682615
rect 244556 679244 244608 679250
rect 244556 679186 244608 679192
rect 244464 450288 244516 450294
rect 244464 450230 244516 450236
rect 244568 449970 244596 679186
rect 245672 461650 245700 684014
rect 247040 683868 247092 683874
rect 247040 683810 247092 683816
rect 245844 680876 245896 680882
rect 245844 680818 245896 680824
rect 245752 680468 245804 680474
rect 245752 680410 245804 680416
rect 245660 461644 245712 461650
rect 245660 461586 245712 461592
rect 244648 456544 244700 456550
rect 244648 456486 244700 456492
rect 241716 449942 241914 449970
rect 241992 449942 242282 449970
rect 242360 449942 242650 449970
rect 242912 449942 243018 449970
rect 243096 449942 243386 449970
rect 243464 449942 243754 449970
rect 243832 449942 244122 449970
rect 244490 449942 244596 449970
rect 244660 449970 244688 456486
rect 244924 456000 244976 456006
rect 244924 455942 244976 455948
rect 244936 449970 244964 455942
rect 245292 450288 245344 450294
rect 245292 450230 245344 450236
rect 245304 449970 245332 450230
rect 245764 449970 245792 680410
rect 245856 466454 245884 680818
rect 245856 466426 246068 466454
rect 246040 449970 246068 466426
rect 246396 461644 246448 461650
rect 246396 461586 246448 461592
rect 246408 449970 246436 461586
rect 244660 449942 244858 449970
rect 244936 449942 245226 449970
rect 245304 449942 245594 449970
rect 245764 449942 245962 449970
rect 246040 449942 246330 449970
rect 246408 449942 246698 449970
rect 247052 449956 247080 683810
rect 247314 682408 247370 682417
rect 247314 682343 247370 682352
rect 247130 682272 247186 682281
rect 247130 682207 247186 682216
rect 247144 449970 247172 682207
rect 247224 681828 247276 681834
rect 247224 681770 247276 681776
rect 247236 456006 247264 681770
rect 247328 466454 247356 682343
rect 247328 466426 247540 466454
rect 247224 456000 247276 456006
rect 247224 455942 247276 455948
rect 247512 449970 247540 466426
rect 247868 456000 247920 456006
rect 247868 455942 247920 455948
rect 247880 449970 247908 455942
rect 248432 449970 248460 684830
rect 248512 683936 248564 683942
rect 248512 683878 248564 683884
rect 248524 450378 248552 683878
rect 248696 681148 248748 681154
rect 248696 681090 248748 681096
rect 248604 680536 248656 680542
rect 248604 680478 248656 680484
rect 248616 451274 248644 680478
rect 248708 466454 248736 681090
rect 248708 466426 249380 466454
rect 248616 451246 249012 451274
rect 248524 450350 248644 450378
rect 248616 449970 248644 450350
rect 248984 449970 249012 451246
rect 249352 449970 249380 466426
rect 249812 450294 249840 684898
rect 252560 684616 252612 684622
rect 252560 684558 252612 684564
rect 249892 681896 249944 681902
rect 249892 681838 249944 681844
rect 249800 450288 249852 450294
rect 249800 450230 249852 450236
rect 249904 449970 249932 681838
rect 249984 681216 250036 681222
rect 249984 681158 250036 681164
rect 249996 451274 250024 681158
rect 251180 681080 251232 681086
rect 251180 681022 251232 681028
rect 250074 679824 250130 679833
rect 250074 679759 250130 679768
rect 250088 466454 250116 679759
rect 250088 466426 250852 466454
rect 249996 451246 250484 451274
rect 250076 450288 250128 450294
rect 250076 450230 250128 450236
rect 250088 449970 250116 450230
rect 250456 449970 250484 451246
rect 250824 449970 250852 466426
rect 251192 456006 251220 681022
rect 251546 462904 251602 462913
rect 251546 462839 251602 462848
rect 251364 459060 251416 459066
rect 251364 459002 251416 459008
rect 251180 456000 251232 456006
rect 251180 455942 251232 455948
rect 251376 449970 251404 459002
rect 251560 449970 251588 462839
rect 251916 456000 251968 456006
rect 251916 455942 251968 455948
rect 251928 449970 251956 455942
rect 252572 450294 252600 684558
rect 252652 683392 252704 683398
rect 252652 683334 252704 683340
rect 252664 456006 252692 683334
rect 252744 682644 252796 682650
rect 252744 682586 252796 682592
rect 252756 458946 252784 682586
rect 260840 682304 260892 682310
rect 260840 682246 260892 682252
rect 259736 682236 259788 682242
rect 259736 682178 259788 682184
rect 256700 682168 256752 682174
rect 256700 682110 256752 682116
rect 255320 682032 255372 682038
rect 255320 681974 255372 681980
rect 254216 681012 254268 681018
rect 254216 680954 254268 680960
rect 252836 680604 252888 680610
rect 252836 680546 252888 680552
rect 252848 463694 252876 680546
rect 254032 679312 254084 679318
rect 254032 679254 254084 679260
rect 252848 463666 253060 463694
rect 252756 458918 252968 458946
rect 252836 458788 252888 458794
rect 252836 458730 252888 458736
rect 252652 456000 252704 456006
rect 252652 455942 252704 455948
rect 252560 450288 252612 450294
rect 252560 450230 252612 450236
rect 247144 449942 247434 449970
rect 247512 449942 247802 449970
rect 247880 449942 248170 449970
rect 248432 449942 248538 449970
rect 248616 449942 248906 449970
rect 248984 449942 249274 449970
rect 249352 449942 249642 449970
rect 249904 449942 250010 449970
rect 250088 449942 250378 449970
rect 250456 449942 250746 449970
rect 250824 449942 251114 449970
rect 251376 449942 251482 449970
rect 251560 449942 251850 449970
rect 251928 449942 252218 449970
rect 232318 449919 232374 449928
rect 193140 449806 193260 449834
rect 193864 449880 193916 449886
rect 193864 449822 193916 449828
rect 193956 449880 194008 449886
rect 193956 449822 194008 449828
rect 201224 449880 201276 449886
rect 201224 449822 201276 449828
rect 229742 449848 229798 449857
rect 193140 449682 193168 449806
rect 193128 449676 193180 449682
rect 193128 449618 193180 449624
rect 193220 449676 193272 449682
rect 193220 449618 193272 449624
rect 193232 449585 193260 449618
rect 193968 449585 193996 449822
rect 200856 449744 200908 449750
rect 195348 449682 195546 449698
rect 200856 449686 200908 449692
rect 195336 449676 195546 449682
rect 195388 449670 195546 449676
rect 195336 449618 195388 449624
rect 200868 449614 200896 449686
rect 201236 449614 201264 449822
rect 252848 449834 252876 458730
rect 252940 451274 252968 458918
rect 253032 458794 253060 463666
rect 253020 458788 253072 458794
rect 253020 458730 253072 458736
rect 253388 456000 253440 456006
rect 253388 455942 253440 455948
rect 252940 451246 253060 451274
rect 252928 450288 252980 450294
rect 252928 450230 252980 450236
rect 252940 449956 252968 450230
rect 253032 449970 253060 451246
rect 253400 449970 253428 455942
rect 253940 451580 253992 451586
rect 253940 451522 253992 451528
rect 253952 449970 253980 451522
rect 254044 450276 254072 679254
rect 254122 678192 254178 678201
rect 254122 678127 254178 678136
rect 254136 453014 254164 678127
rect 254124 453008 254176 453014
rect 254124 452950 254176 452956
rect 254228 451586 254256 680954
rect 254492 460284 254544 460290
rect 254492 460226 254544 460232
rect 254216 451580 254268 451586
rect 254216 451522 254268 451528
rect 254044 450248 254164 450276
rect 254136 449970 254164 450248
rect 254504 449970 254532 460226
rect 255332 453014 255360 681974
rect 255412 680672 255464 680678
rect 255412 680614 255464 680620
rect 254860 453008 254912 453014
rect 254860 452950 254912 452956
rect 255320 453008 255372 453014
rect 255320 452950 255372 452956
rect 254872 449970 254900 452950
rect 255424 449970 255452 680614
rect 255502 679688 255558 679697
rect 255502 679623 255558 679632
rect 255516 460934 255544 679623
rect 255516 460906 256372 460934
rect 255594 457464 255650 457473
rect 255594 457399 255650 457408
rect 255608 449970 255636 457399
rect 255964 453008 256016 453014
rect 255964 452950 256016 452956
rect 255976 449970 256004 452950
rect 256344 449970 256372 460906
rect 256712 452946 256740 682110
rect 258356 682100 258408 682106
rect 258356 682042 258408 682048
rect 256792 681284 256844 681290
rect 256792 681226 256844 681232
rect 256804 453014 256832 681226
rect 256884 680740 256936 680746
rect 256884 680682 256936 680688
rect 256792 453008 256844 453014
rect 256792 452950 256844 452956
rect 256700 452940 256752 452946
rect 256700 452882 256752 452888
rect 256896 449970 256924 680682
rect 258172 679720 258224 679726
rect 258172 679662 258224 679668
rect 258080 458992 258132 458998
rect 258080 458934 258132 458940
rect 258092 453014 258120 458934
rect 257068 453008 257120 453014
rect 257068 452950 257120 452956
rect 258080 453008 258132 453014
rect 258080 452950 258132 452956
rect 257080 449970 257108 452950
rect 257436 452940 257488 452946
rect 257436 452882 257488 452888
rect 257448 449970 257476 452882
rect 258184 449970 258212 679662
rect 258264 679652 258316 679658
rect 258264 679594 258316 679600
rect 258276 453558 258304 679594
rect 258368 460934 258396 682042
rect 259552 681964 259604 681970
rect 259552 681906 259604 681912
rect 258368 460906 258580 460934
rect 258264 453552 258316 453558
rect 258264 453494 258316 453500
rect 258264 453008 258316 453014
rect 258264 452950 258316 452956
rect 253032 449942 253322 449970
rect 253400 449942 253690 449970
rect 253952 449942 254058 449970
rect 254136 449942 254426 449970
rect 254504 449942 254794 449970
rect 254872 449942 255162 449970
rect 255424 449942 255530 449970
rect 255608 449942 255898 449970
rect 255976 449942 256266 449970
rect 256344 449942 256634 449970
rect 256896 449942 257002 449970
rect 257080 449942 257370 449970
rect 257448 449942 257738 449970
rect 258106 449942 258212 449970
rect 258276 449970 258304 452950
rect 258552 449970 258580 460906
rect 259460 458856 259512 458862
rect 259460 458798 259512 458804
rect 258908 453552 258960 453558
rect 258908 453494 258960 453500
rect 258920 449970 258948 453494
rect 259472 449970 259500 458798
rect 259564 453014 259592 681906
rect 259644 679040 259696 679046
rect 259644 678982 259696 678988
rect 259552 453008 259604 453014
rect 259552 452950 259604 452956
rect 259656 452946 259684 678982
rect 259748 456794 259776 682178
rect 259748 456766 259868 456794
rect 259644 452940 259696 452946
rect 259644 452882 259696 452888
rect 259840 449970 259868 456766
rect 260380 453008 260432 453014
rect 260380 452950 260432 452956
rect 260012 452940 260064 452946
rect 260012 452882 260064 452888
rect 260024 449970 260052 452882
rect 260392 449970 260420 452950
rect 260852 449970 260880 682246
rect 262220 497140 262272 497146
rect 262220 497082 262272 497088
rect 260932 497072 260984 497078
rect 260932 497014 260984 497020
rect 260944 453014 260972 497014
rect 261024 467220 261076 467226
rect 261024 467162 261076 467168
rect 261036 456794 261064 467162
rect 261116 463004 261168 463010
rect 261116 462946 261168 462952
rect 261128 460934 261156 462946
rect 261128 460906 261892 460934
rect 261036 456766 261156 456794
rect 260932 453008 260984 453014
rect 260932 452950 260984 452956
rect 261128 449970 261156 456766
rect 261484 453008 261536 453014
rect 261484 452950 261536 452956
rect 261496 449970 261524 452950
rect 261864 449970 261892 460906
rect 262232 453014 262260 497082
rect 262312 494760 262364 494766
rect 262312 494702 262364 494708
rect 262220 453008 262272 453014
rect 262220 452950 262272 452956
rect 262324 449970 262352 494702
rect 262404 487824 262456 487830
rect 262404 487766 262456 487772
rect 262416 460934 262444 487766
rect 263600 483676 263652 483682
rect 263600 483618 263652 483624
rect 262416 460906 262628 460934
rect 262600 449970 262628 460906
rect 263612 453014 263640 483618
rect 266372 476882 266400 697546
rect 271144 696992 271196 696998
rect 271144 696934 271196 696940
rect 270500 535492 270552 535498
rect 270500 535434 270552 535440
rect 269120 496188 269172 496194
rect 269120 496130 269172 496136
rect 266452 486464 266504 486470
rect 266452 486406 266504 486412
rect 266360 476876 266412 476882
rect 266360 476818 266412 476824
rect 266360 475380 266412 475386
rect 266360 475322 266412 475328
rect 264980 474088 265032 474094
rect 264980 474030 265032 474036
rect 263692 472660 263744 472666
rect 263692 472602 263744 472608
rect 262956 453008 263008 453014
rect 262956 452950 263008 452956
rect 263600 453008 263652 453014
rect 263600 452950 263652 452956
rect 262968 449970 262996 452950
rect 263704 449970 263732 472602
rect 263784 461644 263836 461650
rect 263784 461586 263836 461592
rect 263796 460934 263824 461586
rect 263796 460906 264100 460934
rect 263784 453008 263836 453014
rect 263784 452950 263836 452956
rect 258276 449942 258474 449970
rect 258552 449942 258842 449970
rect 258920 449942 259210 449970
rect 259472 449942 259578 449970
rect 259840 449942 259946 449970
rect 260024 449942 260314 449970
rect 260392 449942 260682 449970
rect 260852 449942 261050 449970
rect 261128 449942 261418 449970
rect 261496 449942 261786 449970
rect 261864 449942 262154 449970
rect 262324 449942 262522 449970
rect 262600 449942 262890 449970
rect 262968 449942 263258 449970
rect 263626 449942 263732 449970
rect 263796 449970 263824 452950
rect 264072 449970 264100 460906
rect 264428 460488 264480 460494
rect 264428 460430 264480 460436
rect 264440 449970 264468 460430
rect 264992 449970 265020 474030
rect 265072 461712 265124 461718
rect 265072 461654 265124 461660
rect 265084 460934 265112 461654
rect 265084 460906 265940 460934
rect 265532 458856 265584 458862
rect 265532 458798 265584 458804
rect 265256 457496 265308 457502
rect 265256 457438 265308 457444
rect 265268 449970 265296 457438
rect 265544 449970 265572 458798
rect 265912 449970 265940 460906
rect 266372 449970 266400 475322
rect 266464 450106 266492 486406
rect 267740 476808 267792 476814
rect 267740 476750 267792 476756
rect 266544 464364 266596 464370
rect 266544 464306 266596 464312
rect 266556 456794 266584 464306
rect 266636 463276 266688 463282
rect 266636 463218 266688 463224
rect 266648 460934 266676 463218
rect 266648 460906 267412 460934
rect 266556 456766 267044 456794
rect 266464 450078 266676 450106
rect 266648 449970 266676 450078
rect 267016 449970 267044 456766
rect 267384 449970 267412 460906
rect 267752 449970 267780 476750
rect 267832 468580 267884 468586
rect 267832 468522 267884 468528
rect 267844 456794 267872 468522
rect 267924 464432 267976 464438
rect 267924 464374 267976 464380
rect 267936 460934 267964 464374
rect 267936 460906 268516 460934
rect 267844 456766 268148 456794
rect 268120 449970 268148 456766
rect 268488 449970 268516 460906
rect 269132 453014 269160 496130
rect 269212 479596 269264 479602
rect 269212 479538 269264 479544
rect 269120 453008 269172 453014
rect 269120 452950 269172 452956
rect 269224 449970 269252 479538
rect 269304 478168 269356 478174
rect 269304 478110 269356 478116
rect 269316 453558 269344 478110
rect 269396 465860 269448 465866
rect 269396 465802 269448 465808
rect 269408 460934 269436 465802
rect 269408 460906 269620 460934
rect 269304 453552 269356 453558
rect 269304 453494 269356 453500
rect 269304 453008 269356 453014
rect 269304 452950 269356 452956
rect 263796 449942 263994 449970
rect 264072 449942 264362 449970
rect 264440 449942 264730 449970
rect 264992 449942 265098 449970
rect 265268 449942 265466 449970
rect 265544 449942 265834 449970
rect 265912 449942 266202 449970
rect 266372 449942 266570 449970
rect 266648 449942 266938 449970
rect 267016 449942 267306 449970
rect 267384 449942 267674 449970
rect 267752 449942 268042 449970
rect 268120 449942 268410 449970
rect 268488 449942 268778 449970
rect 269146 449942 269252 449970
rect 269316 449970 269344 452950
rect 269592 449970 269620 460906
rect 269948 453552 270000 453558
rect 269948 453494 270000 453500
rect 269960 449970 269988 453494
rect 270512 450022 270540 535434
rect 270592 481024 270644 481030
rect 270592 480966 270644 480972
rect 270604 452946 270632 480966
rect 271156 478242 271184 696934
rect 280804 532772 280856 532778
rect 280804 532714 280856 532720
rect 279424 529984 279476 529990
rect 279424 529926 279476 529932
rect 277584 509312 277636 509318
rect 277584 509254 277636 509260
rect 276020 497276 276072 497282
rect 276020 497218 276072 497224
rect 271880 496936 271932 496942
rect 271880 496878 271932 496884
rect 271144 478236 271196 478242
rect 271144 478178 271196 478184
rect 270684 471300 270736 471306
rect 270684 471242 270736 471248
rect 270696 453014 270724 471242
rect 270776 469940 270828 469946
rect 270776 469882 270828 469888
rect 270684 453008 270736 453014
rect 270684 452950 270736 452956
rect 270592 452940 270644 452946
rect 270592 452882 270644 452888
rect 270788 452826 270816 469882
rect 271892 453014 271920 496878
rect 274640 496120 274692 496126
rect 274640 496062 274692 496068
rect 273260 493332 273312 493338
rect 273260 493274 273312 493280
rect 271972 482316 272024 482322
rect 271972 482258 272024 482264
rect 271420 453008 271472 453014
rect 271420 452950 271472 452956
rect 271880 453008 271932 453014
rect 271880 452950 271932 452956
rect 271052 452940 271104 452946
rect 271052 452882 271104 452888
rect 270604 452798 270816 452826
rect 270500 450016 270552 450022
rect 269316 449942 269514 449970
rect 269592 449942 269882 449970
rect 269960 449942 270250 449970
rect 270500 449958 270552 449964
rect 270604 449956 270632 452798
rect 270776 450016 270828 450022
rect 271064 449970 271092 452882
rect 271432 449970 271460 452950
rect 271984 449970 272012 482258
rect 272156 460284 272208 460290
rect 272156 460226 272208 460232
rect 272168 449970 272196 460226
rect 273272 455818 273300 493274
rect 273352 469872 273404 469878
rect 273352 469814 273404 469820
rect 273364 456006 273392 469814
rect 273444 468512 273496 468518
rect 273444 468454 273496 468460
rect 273456 460934 273484 468454
rect 273456 460906 273668 460934
rect 273352 456000 273404 456006
rect 273352 455942 273404 455948
rect 273272 455790 273576 455818
rect 273444 455660 273496 455666
rect 273444 455602 273496 455608
rect 273168 453552 273220 453558
rect 273168 453494 273220 453500
rect 272524 453008 272576 453014
rect 272524 452950 272576 452956
rect 272536 449970 272564 452950
rect 270828 449964 270986 449970
rect 270776 449958 270986 449964
rect 270788 449942 270986 449958
rect 271064 449942 271354 449970
rect 271432 449942 271722 449970
rect 271984 449942 272090 449970
rect 272168 449942 272458 449970
rect 272536 449942 272826 449970
rect 273180 449956 273208 453494
rect 273456 449970 273484 455602
rect 273548 451274 273576 455790
rect 273640 455666 273668 460906
rect 273996 456000 274048 456006
rect 273996 455942 274048 455948
rect 273628 455660 273680 455666
rect 273628 455602 273680 455608
rect 273548 451246 273668 451274
rect 273640 449970 273668 451246
rect 274008 449970 274036 455942
rect 273456 449942 273562 449970
rect 273640 449942 273930 449970
rect 274008 449942 274298 449970
rect 274652 449956 274680 496062
rect 274732 490612 274784 490618
rect 274732 490554 274784 490560
rect 274744 450294 274772 490554
rect 274824 465792 274876 465798
rect 274824 465734 274876 465740
rect 274836 460934 274864 465734
rect 274836 460906 274956 460934
rect 274732 450288 274784 450294
rect 274732 450230 274784 450236
rect 274928 449970 274956 460906
rect 275468 460216 275520 460222
rect 275468 460158 275520 460164
rect 275100 450288 275152 450294
rect 275100 450230 275152 450236
rect 275112 449970 275140 450230
rect 275480 449970 275508 460158
rect 276032 456278 276060 497218
rect 277492 497004 277544 497010
rect 277492 496946 277544 496952
rect 276112 491972 276164 491978
rect 276112 491914 276164 491920
rect 276020 456272 276072 456278
rect 276020 456214 276072 456220
rect 276124 456006 276152 491914
rect 276204 489252 276256 489258
rect 276204 489194 276256 489200
rect 276112 456000 276164 456006
rect 276112 455942 276164 455948
rect 276216 449970 276244 489194
rect 276296 467152 276348 467158
rect 276296 467094 276348 467100
rect 274928 449942 275034 449970
rect 275112 449942 275402 449970
rect 275480 449942 275770 449970
rect 276138 449942 276244 449970
rect 276308 449970 276336 467094
rect 276940 456272 276992 456278
rect 276940 456214 276992 456220
rect 276572 456000 276624 456006
rect 276572 455942 276624 455948
rect 276584 449970 276612 455942
rect 276952 449970 276980 456214
rect 277504 449970 277532 496946
rect 277596 460934 277624 509254
rect 279436 463282 279464 529926
rect 280816 465866 280844 532714
rect 282932 492046 282960 702406
rect 295984 527196 296036 527202
rect 295984 527138 296036 527144
rect 283564 497208 283616 497214
rect 283564 497150 283616 497156
rect 282920 492040 282972 492046
rect 282920 491982 282972 491988
rect 280804 465860 280856 465866
rect 280804 465802 280856 465808
rect 279424 463276 279476 463282
rect 279424 463218 279476 463224
rect 277596 460906 277716 460934
rect 277688 449970 277716 460906
rect 280988 460556 281040 460562
rect 280988 460498 281040 460504
rect 280250 458960 280306 458969
rect 280250 458895 280306 458904
rect 278688 457224 278740 457230
rect 278688 457166 278740 457172
rect 278700 454986 278728 457166
rect 279516 456204 279568 456210
rect 279516 456146 279568 456152
rect 278044 454980 278096 454986
rect 278044 454922 278096 454928
rect 278688 454980 278740 454986
rect 278688 454922 278740 454928
rect 278056 449970 278084 454922
rect 278780 451308 278832 451314
rect 278780 451250 278832 451256
rect 278792 450566 278820 451250
rect 279424 451036 279476 451042
rect 279424 450978 279476 450984
rect 278780 450560 278832 450566
rect 278780 450502 278832 450508
rect 279054 449984 279110 449993
rect 276308 449942 276506 449970
rect 276584 449942 276874 449970
rect 276952 449942 277242 449970
rect 277504 449942 277610 449970
rect 277688 449942 277978 449970
rect 278056 449942 278346 449970
rect 278516 449954 278714 449970
rect 278504 449948 278714 449954
rect 278556 449942 278714 449948
rect 279436 449956 279464 450978
rect 279528 449970 279556 456146
rect 280158 451752 280214 451761
rect 280158 451687 280214 451696
rect 279528 449942 279818 449970
rect 280172 449956 280200 451687
rect 280264 449970 280292 458895
rect 280896 450968 280948 450974
rect 280896 450910 280948 450916
rect 280264 449942 280554 449970
rect 280908 449956 280936 450910
rect 281000 449970 281028 460498
rect 282184 456272 282236 456278
rect 282184 456214 282236 456220
rect 282196 451518 282224 456214
rect 282460 456204 282512 456210
rect 282460 456146 282512 456152
rect 282472 453490 282500 456146
rect 283010 455696 283066 455705
rect 283010 455631 283066 455640
rect 282460 453484 282512 453490
rect 282460 453426 282512 453432
rect 282368 451784 282420 451790
rect 282368 451726 282420 451732
rect 282380 451586 282408 451726
rect 282368 451580 282420 451586
rect 282368 451522 282420 451528
rect 282184 451512 282236 451518
rect 282184 451454 282236 451460
rect 281632 450832 281684 450838
rect 281632 450774 281684 450780
rect 281000 449942 281290 449970
rect 281644 449956 281672 450774
rect 282196 449970 282224 451454
rect 282026 449942 282224 449970
rect 282380 449956 282408 451522
rect 282472 449970 282500 453426
rect 283024 449970 283052 455631
rect 283194 454608 283250 454617
rect 283194 454543 283250 454552
rect 283208 449970 283236 454543
rect 283576 453558 283604 497150
rect 294144 463208 294196 463214
rect 294144 463150 294196 463156
rect 288714 462632 288770 462641
rect 288714 462567 288770 462576
rect 284298 462496 284354 462505
rect 284298 462431 284354 462440
rect 284312 460934 284340 462431
rect 288728 460934 288756 462567
rect 290004 461780 290056 461786
rect 290004 461722 290056 461728
rect 284312 460906 284708 460934
rect 288728 460906 289124 460934
rect 283656 459128 283708 459134
rect 283656 459070 283708 459076
rect 283564 453552 283616 453558
rect 283564 453494 283616 453500
rect 283668 451274 283696 459070
rect 283930 454064 283986 454073
rect 283930 453999 283986 454008
rect 283576 451246 283696 451274
rect 283576 449970 283604 451246
rect 283944 449970 283972 453999
rect 284576 450764 284628 450770
rect 284576 450706 284628 450712
rect 282472 449942 282762 449970
rect 283024 449942 283130 449970
rect 283208 449942 283498 449970
rect 283576 449942 283866 449970
rect 283944 449942 284234 449970
rect 284588 449956 284616 450706
rect 284680 449970 284708 460906
rect 286508 459808 286560 459814
rect 286508 459750 286560 459756
rect 285862 456104 285918 456113
rect 285862 456039 285918 456048
rect 285036 454436 285088 454442
rect 285036 454378 285088 454384
rect 285048 449970 285076 454378
rect 285876 449970 285904 456039
rect 285956 454912 286008 454918
rect 285956 454854 286008 454860
rect 284680 449942 284970 449970
rect 285048 449942 285338 449970
rect 285706 449942 285904 449970
rect 285968 449970 285996 454854
rect 286520 452130 286548 459750
rect 287980 458788 288032 458794
rect 287980 458730 288032 458736
rect 287610 457328 287666 457337
rect 287610 457263 287666 457272
rect 287152 452940 287204 452946
rect 287152 452882 287204 452888
rect 286508 452124 286560 452130
rect 286508 452066 286560 452072
rect 286416 451716 286468 451722
rect 286416 451658 286468 451664
rect 285968 449942 286074 449970
rect 286428 449956 286456 451658
rect 286520 449970 286548 452066
rect 286520 449942 286810 449970
rect 287164 449956 287192 452882
rect 287520 452736 287572 452742
rect 287520 452678 287572 452684
rect 287532 449956 287560 452678
rect 287624 449970 287652 457263
rect 287992 449970 288020 458730
rect 288440 457632 288492 457638
rect 288440 457574 288492 457580
rect 288452 449970 288480 457574
rect 288716 456884 288768 456890
rect 288716 456826 288768 456832
rect 288728 449970 288756 456826
rect 289096 449970 289124 460906
rect 289268 457632 289320 457638
rect 289268 457574 289320 457580
rect 289280 457201 289308 457574
rect 289266 457192 289322 457201
rect 289266 457127 289322 457136
rect 289452 454368 289504 454374
rect 289452 454310 289504 454316
rect 289464 449970 289492 454310
rect 290016 449970 290044 461722
rect 294156 460934 294184 463150
rect 294156 460906 294276 460934
rect 292764 459876 292816 459882
rect 292764 459818 292816 459824
rect 291200 458448 291252 458454
rect 291200 458390 291252 458396
rect 291212 452130 291240 458390
rect 292026 457464 292082 457473
rect 292026 457399 292082 457408
rect 291660 453620 291712 453626
rect 291660 453562 291712 453568
rect 291672 453014 291700 453562
rect 291934 453520 291990 453529
rect 291934 453455 291990 453464
rect 291660 453008 291712 453014
rect 291660 452950 291712 452956
rect 291200 452124 291252 452130
rect 291200 452066 291252 452072
rect 290464 452056 290516 452062
rect 290464 451998 290516 452004
rect 287624 449942 287914 449970
rect 287992 449942 288282 449970
rect 288452 449942 288650 449970
rect 288728 449942 289018 449970
rect 289096 449942 289386 449970
rect 289464 449942 289754 449970
rect 290016 449942 290122 449970
rect 290476 449956 290504 451998
rect 290832 451512 290884 451518
rect 290832 451454 290884 451460
rect 290556 450084 290608 450090
rect 290556 450026 290608 450032
rect 290568 449970 290596 450026
rect 290844 449970 290872 451454
rect 290568 449956 290872 449970
rect 291212 449956 291240 452066
rect 291672 449970 291700 452950
rect 290568 449942 290858 449956
rect 291594 449942 291700 449970
rect 291948 449956 291976 453455
rect 292040 449970 292068 457399
rect 292776 449970 292804 459818
rect 292856 457564 292908 457570
rect 292856 457506 292908 457512
rect 292040 449942 292330 449970
rect 292698 449942 292804 449970
rect 292868 449970 292896 457506
rect 293408 456340 293460 456346
rect 293408 456282 293460 456288
rect 292868 449942 293066 449970
rect 293420 449956 293448 456282
rect 294144 454300 294196 454306
rect 294144 454242 294196 454248
rect 293776 450560 293828 450566
rect 293776 450502 293828 450508
rect 293788 449956 293816 450502
rect 294156 449956 294184 454242
rect 294248 449970 294276 460906
rect 295996 460494 296024 527138
rect 298744 507884 298796 507890
rect 298744 507826 298796 507832
rect 298756 467226 298784 507826
rect 299492 472734 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 331232 504422 331260 702986
rect 348804 699718 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 345664 699712 345716 699718
rect 345664 699654 345716 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 345676 507142 345704 699654
rect 345664 507136 345716 507142
rect 345664 507078 345716 507084
rect 331220 504416 331272 504422
rect 331220 504358 331272 504364
rect 364352 502994 364380 702406
rect 371884 700392 371936 700398
rect 371884 700334 371936 700340
rect 371896 505782 371924 700334
rect 397472 699718 397500 703520
rect 413664 700330 413692 703520
rect 429856 700330 429884 703520
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 418804 700324 418856 700330
rect 418804 700266 418856 700272
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 390650 682544 390706 682553
rect 390650 682479 390706 682488
rect 390558 682000 390614 682009
rect 390558 681935 390614 681944
rect 389178 679008 389234 679017
rect 389178 678943 389234 678952
rect 371884 505776 371936 505782
rect 371884 505718 371936 505724
rect 364340 502988 364392 502994
rect 364340 502930 364392 502936
rect 299480 472728 299532 472734
rect 299480 472670 299532 472676
rect 298744 467220 298796 467226
rect 298744 467162 298796 467168
rect 367100 465520 367152 465526
rect 367100 465462 367152 465468
rect 327356 464636 327408 464642
rect 327356 464578 327408 464584
rect 316316 464568 316368 464574
rect 316316 464510 316368 464516
rect 302240 464500 302292 464506
rect 302240 464442 302292 464448
rect 298192 463140 298244 463146
rect 298192 463082 298244 463088
rect 295984 460488 296036 460494
rect 295984 460430 296036 460436
rect 297548 460420 297600 460426
rect 297548 460362 297600 460368
rect 296812 458720 296864 458726
rect 296812 458662 296864 458668
rect 296718 457192 296774 457201
rect 296718 457127 296774 457136
rect 295984 455048 296036 455054
rect 295984 454990 296036 454996
rect 295996 453490 296024 454990
rect 295984 453484 296036 453490
rect 295984 453426 296036 453432
rect 294880 452260 294932 452266
rect 294880 452202 294932 452208
rect 294248 449942 294538 449970
rect 294892 449956 294920 452202
rect 295246 452024 295302 452033
rect 295246 451959 295302 451968
rect 295616 451988 295668 451994
rect 295260 450702 295288 451959
rect 295616 451930 295668 451936
rect 295248 450696 295300 450702
rect 295248 450638 295300 450644
rect 295260 449956 295288 450638
rect 295628 449956 295656 451930
rect 295996 449956 296024 453426
rect 296352 451308 296404 451314
rect 296352 451250 296404 451256
rect 296364 449956 296392 451250
rect 296732 449956 296760 457127
rect 296824 449970 296852 458662
rect 297180 457428 297232 457434
rect 297180 457370 297232 457376
rect 297192 449970 297220 457370
rect 297364 452124 297416 452130
rect 297364 452066 297416 452072
rect 297376 451790 297404 452066
rect 297364 451784 297416 451790
rect 297364 451726 297416 451732
rect 297560 449970 297588 460362
rect 297640 451988 297692 451994
rect 297640 451930 297692 451936
rect 297652 451874 297680 451930
rect 297824 451920 297876 451926
rect 297652 451868 297824 451874
rect 297652 451862 297876 451868
rect 297652 451846 297864 451862
rect 298204 450770 298232 463082
rect 298284 462392 298336 462398
rect 298284 462334 298336 462340
rect 298192 450764 298244 450770
rect 298192 450706 298244 450712
rect 298296 449970 298324 462334
rect 301596 460352 301648 460358
rect 301596 460294 301648 460300
rect 301044 460148 301096 460154
rect 301044 460090 301096 460096
rect 299664 458924 299716 458930
rect 299664 458866 299716 458872
rect 299480 455116 299532 455122
rect 299480 455058 299532 455064
rect 299492 453558 299520 455058
rect 299480 453552 299532 453558
rect 299480 453494 299532 453500
rect 299676 452538 299704 458866
rect 300490 457600 300546 457609
rect 300490 457535 300546 457544
rect 300032 453552 300084 453558
rect 300032 453494 300084 453500
rect 299664 452532 299716 452538
rect 299664 452474 299716 452480
rect 299296 451444 299348 451450
rect 299296 451386 299348 451392
rect 298652 450764 298704 450770
rect 298652 450706 298704 450712
rect 298560 450696 298612 450702
rect 298560 450638 298612 450644
rect 296824 449942 297114 449970
rect 297192 449942 297482 449970
rect 297560 449942 297850 449970
rect 298218 449942 298324 449970
rect 298572 449956 298600 450638
rect 298664 449970 298692 450706
rect 298664 449942 298954 449970
rect 299308 449956 299336 451386
rect 299676 449956 299704 452474
rect 300044 449956 300072 453494
rect 300398 453384 300454 453393
rect 300398 453319 300454 453328
rect 300412 449956 300440 453319
rect 300504 449970 300532 457535
rect 301056 449970 301084 460090
rect 301228 457360 301280 457366
rect 301228 457302 301280 457308
rect 301240 449970 301268 457302
rect 301608 449970 301636 460294
rect 302252 450294 302280 464442
rect 302332 463072 302384 463078
rect 302332 463014 302384 463020
rect 302344 453082 302372 463014
rect 306380 462936 306432 462942
rect 306380 462878 306432 462884
rect 302422 462768 302478 462777
rect 302422 462703 302478 462712
rect 302436 456794 302464 462703
rect 305000 462460 305052 462466
rect 305000 462402 305052 462408
rect 305012 460934 305040 462402
rect 306392 460934 306420 462878
rect 309140 462868 309192 462874
rect 309140 462810 309192 462816
rect 309152 460934 309180 462810
rect 314660 462800 314712 462806
rect 314660 462742 314712 462748
rect 310520 462664 310572 462670
rect 310520 462606 310572 462612
rect 310532 460934 310560 462606
rect 313280 461780 313332 461786
rect 313280 461722 313332 461728
rect 313292 460934 313320 461722
rect 305012 460906 306052 460934
rect 306392 460906 306788 460934
rect 309152 460906 310100 460934
rect 310532 460906 310652 460934
rect 313292 460906 313780 460934
rect 305644 459944 305696 459950
rect 305644 459886 305696 459892
rect 305184 458924 305236 458930
rect 305184 458866 305236 458872
rect 303988 458312 304040 458318
rect 303988 458254 304040 458260
rect 302436 456766 302556 456794
rect 302332 453076 302384 453082
rect 302332 453018 302384 453024
rect 302528 450650 302556 456766
rect 302700 453076 302752 453082
rect 302700 453018 302752 453024
rect 302344 450622 302556 450650
rect 302240 450288 302292 450294
rect 302240 450230 302292 450236
rect 302344 449970 302372 450622
rect 302424 450288 302476 450294
rect 302424 450230 302476 450236
rect 300504 449942 300794 449970
rect 301056 449942 301162 449970
rect 301240 449942 301530 449970
rect 301608 449942 301898 449970
rect 302266 449942 302372 449970
rect 302436 449970 302464 450230
rect 302712 449970 302740 453018
rect 303896 452532 303948 452538
rect 303896 452474 303948 452480
rect 303712 452192 303764 452198
rect 303712 452134 303764 452140
rect 303724 451926 303752 452134
rect 303908 452062 303936 452474
rect 304000 452130 304028 458254
rect 304814 455696 304870 455705
rect 304814 455631 304870 455640
rect 304080 454232 304132 454238
rect 304080 454174 304132 454180
rect 304724 454232 304776 454238
rect 304724 454174 304776 454180
rect 303988 452124 304040 452130
rect 303988 452066 304040 452072
rect 303896 452056 303948 452062
rect 303896 451998 303948 452004
rect 303712 451920 303764 451926
rect 303712 451862 303764 451868
rect 303342 451616 303398 451625
rect 303342 451551 303398 451560
rect 302436 449942 302634 449970
rect 302712 449942 303002 449970
rect 303356 449956 303384 451551
rect 304000 449970 304028 452066
rect 303738 449942 304028 449970
rect 304092 449956 304120 454174
rect 304736 453626 304764 454174
rect 304724 453620 304776 453626
rect 304724 453562 304776 453568
rect 304446 453384 304502 453393
rect 304446 453319 304502 453328
rect 304264 452192 304316 452198
rect 304264 452134 304316 452140
rect 304276 451994 304304 452134
rect 304264 451988 304316 451994
rect 304264 451930 304316 451936
rect 304460 449956 304488 453319
rect 304828 449956 304856 455631
rect 305196 449956 305224 458866
rect 305550 453248 305606 453257
rect 305550 453183 305606 453192
rect 305564 449956 305592 453183
rect 305656 449970 305684 459886
rect 306024 449970 306052 460906
rect 306656 455048 306708 455054
rect 306656 454990 306708 454996
rect 305656 449942 305946 449970
rect 306024 449942 306314 449970
rect 306668 449956 306696 454990
rect 306760 449970 306788 460906
rect 309232 460352 309284 460358
rect 309232 460294 309284 460300
rect 308588 457088 308640 457094
rect 308588 457030 308640 457036
rect 308128 454164 308180 454170
rect 308128 454106 308180 454112
rect 308140 452810 308168 454106
rect 308128 452804 308180 452810
rect 308128 452746 308180 452752
rect 307760 451920 307812 451926
rect 307760 451862 307812 451868
rect 306760 449942 307050 449970
rect 307772 449956 307800 451862
rect 308140 449956 308168 452746
rect 308494 451616 308550 451625
rect 308494 451551 308550 451560
rect 308508 449956 308536 451551
rect 308600 449970 308628 457030
rect 308600 449942 308890 449970
rect 309244 449956 309272 460294
rect 309414 457736 309470 457745
rect 309414 457671 309470 457680
rect 309428 449970 309456 457671
rect 309968 454776 310020 454782
rect 309968 454718 310020 454724
rect 309428 449942 309626 449970
rect 309980 449956 310008 454718
rect 310072 449970 310100 460906
rect 310624 456794 310652 460906
rect 312636 458652 312688 458658
rect 312636 458594 312688 458600
rect 310624 456766 310836 456794
rect 310520 454708 310572 454714
rect 310520 454650 310572 454656
rect 310532 451314 310560 454650
rect 310704 454232 310756 454238
rect 310704 454174 310756 454180
rect 310520 451308 310572 451314
rect 310520 451250 310572 451256
rect 310072 449942 310362 449970
rect 310716 449956 310744 454174
rect 310808 449970 310836 456766
rect 311440 456068 311492 456074
rect 311440 456010 311492 456016
rect 310808 449942 311098 449970
rect 311452 449956 311480 456010
rect 312268 456000 312320 456006
rect 312268 455942 312320 455948
rect 312176 454096 312228 454102
rect 312176 454038 312228 454044
rect 312188 452878 312216 454038
rect 312176 452872 312228 452878
rect 312176 452814 312228 452820
rect 311808 451308 311860 451314
rect 311808 451250 311860 451256
rect 311820 449956 311848 451250
rect 312188 449956 312216 452814
rect 312280 449970 312308 455942
rect 312648 449970 312676 458594
rect 313372 455592 313424 455598
rect 313372 455534 313424 455540
rect 313384 449970 313412 455534
rect 313646 452976 313702 452985
rect 313646 452911 313702 452920
rect 312280 449942 312570 449970
rect 312648 449942 312938 449970
rect 313306 449942 313412 449970
rect 313660 449956 313688 452911
rect 313752 449970 313780 460906
rect 314108 454708 314160 454714
rect 314108 454650 314160 454656
rect 314120 449970 314148 454650
rect 314672 449970 314700 462742
rect 316328 460934 316356 464510
rect 320364 464296 320416 464302
rect 320364 464238 320416 464244
rect 317420 462732 317472 462738
rect 317420 462674 317472 462680
rect 317432 460934 317460 462674
rect 320376 460934 320404 464238
rect 323124 462732 323176 462738
rect 323124 462674 323176 462680
rect 323136 460934 323164 462674
rect 327368 460934 327396 464578
rect 331496 464228 331548 464234
rect 331496 464170 331548 464176
rect 330116 462800 330168 462806
rect 330116 462742 330168 462748
rect 330128 460934 330156 462742
rect 316328 460906 317092 460934
rect 317432 460906 317828 460934
rect 320376 460906 320772 460934
rect 323136 460906 323716 460934
rect 327368 460906 327764 460934
rect 330128 460906 330340 460934
rect 316132 460488 316184 460494
rect 316132 460430 316184 460436
rect 315578 456104 315634 456113
rect 315578 456039 315634 456048
rect 315118 452296 315174 452305
rect 315118 452231 315174 452240
rect 314752 451852 314804 451858
rect 314752 451794 314804 451800
rect 314764 451450 314792 451794
rect 314752 451444 314804 451450
rect 314752 451386 314804 451392
rect 313752 449942 314042 449970
rect 314120 449942 314410 449970
rect 314672 449942 314778 449970
rect 315132 449956 315160 452231
rect 315488 451444 315540 451450
rect 315488 451386 315540 451392
rect 315500 449956 315528 451386
rect 315592 449970 315620 456039
rect 316144 449970 316172 460430
rect 316684 456952 316736 456958
rect 316684 456894 316736 456900
rect 316316 455932 316368 455938
rect 316316 455874 316368 455880
rect 316328 449970 316356 455874
rect 316696 449970 316724 456894
rect 317064 449970 317092 460906
rect 317512 454912 317564 454918
rect 317512 454854 317564 454860
rect 317524 449970 317552 454854
rect 317800 449970 317828 460906
rect 318800 460420 318852 460426
rect 318800 460362 318852 460368
rect 318430 453112 318486 453121
rect 318430 453047 318486 453056
rect 315592 449942 315882 449970
rect 316144 449942 316250 449970
rect 316328 449942 316618 449970
rect 316696 449942 316986 449970
rect 317064 449942 317354 449970
rect 317524 449942 317722 449970
rect 317800 449942 318090 449970
rect 318444 449956 318472 453047
rect 318812 451654 318840 460362
rect 319628 459264 319680 459270
rect 319628 459206 319680 459212
rect 319260 458312 319312 458318
rect 319260 458254 319312 458260
rect 318984 457292 319036 457298
rect 318984 457234 319036 457240
rect 318800 451648 318852 451654
rect 318800 451590 318852 451596
rect 318812 449956 318840 451590
rect 318996 449970 319024 457234
rect 319272 449970 319300 458254
rect 319640 449970 319668 459206
rect 320180 457020 320232 457026
rect 320180 456962 320232 456968
rect 320192 449970 320220 456962
rect 320640 450628 320692 450634
rect 320640 450570 320692 450576
rect 318996 449942 319194 449970
rect 319272 449942 319562 449970
rect 319640 449942 319930 449970
rect 320192 449942 320298 449970
rect 320652 449956 320680 450570
rect 320744 449970 320772 460906
rect 321098 460184 321154 460193
rect 321098 460119 321154 460128
rect 320824 451852 320876 451858
rect 320824 451794 320876 451800
rect 320836 451450 320864 451794
rect 320824 451444 320876 451450
rect 320824 451386 320876 451392
rect 321112 449970 321140 460119
rect 323124 458584 323176 458590
rect 323124 458526 323176 458532
rect 322204 455864 322256 455870
rect 322204 455806 322256 455812
rect 321836 454844 321888 454850
rect 321836 454786 321888 454792
rect 321744 450492 321796 450498
rect 321744 450434 321796 450440
rect 320744 449942 321034 449970
rect 321112 449942 321402 449970
rect 321756 449956 321784 450434
rect 321848 449970 321876 454786
rect 322216 449970 322244 455806
rect 322940 455728 322992 455734
rect 322940 455670 322992 455676
rect 322846 450528 322902 450537
rect 322846 450463 322902 450472
rect 321848 449942 322138 449970
rect 322216 449942 322506 449970
rect 322860 449956 322888 450463
rect 322952 450294 322980 455670
rect 322940 450288 322992 450294
rect 322940 450230 322992 450236
rect 323136 449970 323164 458526
rect 323308 450288 323360 450294
rect 323308 450230 323360 450236
rect 323320 449970 323348 450230
rect 323688 449970 323716 460906
rect 324502 458824 324558 458833
rect 324502 458759 324558 458768
rect 327170 458824 327226 458833
rect 327170 458759 327226 458768
rect 324318 452704 324374 452713
rect 324318 452639 324374 452648
rect 323136 449942 323242 449970
rect 323320 449942 323610 449970
rect 323688 449942 323978 449970
rect 324332 449956 324360 452639
rect 324516 449970 324544 458759
rect 325700 458584 325752 458590
rect 325700 458526 325752 458532
rect 325056 453416 325108 453422
rect 325056 453358 325108 453364
rect 324516 449942 324714 449970
rect 325068 449956 325096 453358
rect 325424 452260 325476 452266
rect 325424 452202 325476 452208
rect 325436 451382 325464 452202
rect 325424 451376 325476 451382
rect 325424 451318 325476 451324
rect 325436 449956 325464 451318
rect 325712 450022 325740 458526
rect 326620 457904 326672 457910
rect 326620 457846 326672 457852
rect 325976 457156 326028 457162
rect 325976 457098 326028 457104
rect 325988 450106 326016 457098
rect 326250 457056 326306 457065
rect 326250 456991 326306 457000
rect 325804 450078 326016 450106
rect 325700 450016 325752 450022
rect 325700 449958 325752 449964
rect 325804 449956 325832 450078
rect 325976 450016 326028 450022
rect 326264 449970 326292 456991
rect 326632 449970 326660 457846
rect 327184 449970 327212 458759
rect 327630 453112 327686 453121
rect 327630 453047 327686 453056
rect 326028 449964 326186 449970
rect 325976 449958 326186 449964
rect 325988 449942 326186 449958
rect 326264 449942 326554 449970
rect 326632 449942 326922 449970
rect 327184 449942 327290 449970
rect 327644 449956 327672 453047
rect 327736 449970 327764 460906
rect 328552 459196 328604 459202
rect 328552 459138 328604 459144
rect 328564 456550 328592 459138
rect 329932 458516 329984 458522
rect 329932 458458 329984 458464
rect 329196 458448 329248 458454
rect 329196 458390 329248 458396
rect 328552 456544 328604 456550
rect 328552 456486 328604 456492
rect 328368 453348 328420 453354
rect 328368 453290 328420 453296
rect 327736 449942 328026 449970
rect 328380 449956 328408 453290
rect 328564 449970 328592 456486
rect 328828 454980 328880 454986
rect 328828 454922 328880 454928
rect 328840 449970 328868 454922
rect 329208 449970 329236 458390
rect 329944 449970 329972 458458
rect 330024 455796 330076 455802
rect 330024 455738 330076 455744
rect 328564 449942 328762 449970
rect 328840 449942 329130 449970
rect 329208 449942 329498 449970
rect 329866 449942 329972 449970
rect 330036 449970 330064 455738
rect 330312 449970 330340 460906
rect 331220 456136 331272 456142
rect 331220 456078 331272 456084
rect 331232 454850 331260 456078
rect 331220 454844 331272 454850
rect 331220 454786 331272 454792
rect 330942 453248 330998 453257
rect 330942 453183 330998 453192
rect 330036 449942 330234 449970
rect 330312 449942 330602 449970
rect 330956 449956 330984 453183
rect 331508 449970 331536 464170
rect 333980 464160 334032 464166
rect 333980 464102 334032 464108
rect 349158 464128 349214 464137
rect 332692 458516 332744 458522
rect 332692 458458 332744 458464
rect 332140 457020 332192 457026
rect 332140 456962 332192 456968
rect 331772 454844 331824 454850
rect 331772 454786 331824 454792
rect 331680 453280 331732 453286
rect 331680 453222 331732 453228
rect 331338 449942 331536 449970
rect 331692 449956 331720 453222
rect 331784 449970 331812 454786
rect 332152 449970 332180 456962
rect 332704 449970 332732 458458
rect 333610 458416 333666 458425
rect 333610 458351 333666 458360
rect 333244 457700 333296 457706
rect 333244 457642 333296 457648
rect 332874 456920 332930 456929
rect 332874 456855 332930 456864
rect 332888 449970 332916 456855
rect 333256 449970 333284 457642
rect 333624 449970 333652 458351
rect 333992 456346 334020 464102
rect 336740 464092 336792 464098
rect 349158 464063 349214 464072
rect 336740 464034 336792 464040
rect 334072 461576 334124 461582
rect 334072 461518 334124 461524
rect 333980 456340 334032 456346
rect 333980 456282 334032 456288
rect 334084 449970 334112 461518
rect 336188 459332 336240 459338
rect 336188 459274 336240 459280
rect 335452 457360 335504 457366
rect 335452 457302 335504 457308
rect 334348 456340 334400 456346
rect 334348 456282 334400 456288
rect 334360 449970 334388 456282
rect 335360 452192 335412 452198
rect 335360 452134 335412 452140
rect 334992 450424 335044 450430
rect 334992 450366 335044 450372
rect 331784 449942 332074 449970
rect 332152 449942 332442 449970
rect 332704 449942 332810 449970
rect 332888 449942 333178 449970
rect 333256 449942 333546 449970
rect 333624 449942 333914 449970
rect 334084 449942 334282 449970
rect 334360 449942 334650 449970
rect 335004 449956 335032 450366
rect 335372 449956 335400 452134
rect 335464 449970 335492 457302
rect 336096 450424 336148 450430
rect 336096 450366 336148 450372
rect 335464 449942 335754 449970
rect 336108 449956 336136 450366
rect 336200 449970 336228 459274
rect 336752 456142 336780 464034
rect 341156 464024 341208 464030
rect 341156 463966 341208 463972
rect 336832 462936 336884 462942
rect 336832 462878 336884 462884
rect 336844 460934 336872 462878
rect 339500 462664 339552 462670
rect 339500 462606 339552 462612
rect 339512 460934 339540 462606
rect 336844 460906 336964 460934
rect 339512 460906 340276 460934
rect 336740 456136 336792 456142
rect 336740 456078 336792 456084
rect 336648 452192 336700 452198
rect 336648 452134 336700 452140
rect 336660 451654 336688 452134
rect 336648 451648 336700 451654
rect 336648 451590 336700 451596
rect 336936 449970 336964 460906
rect 338396 460012 338448 460018
rect 338396 459954 338448 459960
rect 337660 456136 337712 456142
rect 337660 456078 337712 456084
rect 337568 453076 337620 453082
rect 337568 453018 337620 453024
rect 336200 449942 336490 449970
rect 336936 449942 337226 449970
rect 337580 449956 337608 453018
rect 337672 449970 337700 456078
rect 338120 453212 338172 453218
rect 338120 453154 338172 453160
rect 338132 449970 338160 453154
rect 338408 449970 338436 459954
rect 339868 458380 339920 458386
rect 339868 458322 339920 458328
rect 338764 457428 338816 457434
rect 338764 457370 338816 457376
rect 338776 449970 338804 457370
rect 339132 455932 339184 455938
rect 339132 455874 339184 455880
rect 339144 449970 339172 455874
rect 339776 450356 339828 450362
rect 339776 450298 339828 450304
rect 337672 449942 337962 449970
rect 338132 449942 338330 449970
rect 338408 449942 338698 449970
rect 338776 449942 339066 449970
rect 339144 449942 339434 449970
rect 339788 449956 339816 450298
rect 339880 449970 339908 458322
rect 340248 449970 340276 460906
rect 340880 453348 340932 453354
rect 340880 453290 340932 453296
rect 339880 449942 340170 449970
rect 340248 449942 340538 449970
rect 340892 449956 340920 453290
rect 341168 449970 341196 463966
rect 343640 463956 343692 463962
rect 343640 463898 343692 463904
rect 342260 463072 342312 463078
rect 342260 463014 342312 463020
rect 341708 456952 341760 456958
rect 341708 456894 341760 456900
rect 341616 453688 341668 453694
rect 341616 453630 341668 453636
rect 341168 449942 341274 449970
rect 341628 449956 341656 453630
rect 341720 449970 341748 456894
rect 342272 453218 342300 463014
rect 342352 461984 342404 461990
rect 342352 461926 342404 461932
rect 342364 460934 342392 461926
rect 342364 460906 342852 460934
rect 342534 458688 342590 458697
rect 342534 458623 342590 458632
rect 342444 458380 342496 458386
rect 342444 458322 342496 458328
rect 342260 453212 342312 453218
rect 342260 453154 342312 453160
rect 342456 449970 342484 458322
rect 341720 449942 342010 449970
rect 342378 449942 342484 449970
rect 342548 449970 342576 458623
rect 342824 449970 342852 460906
rect 343652 456794 343680 463898
rect 346584 463888 346636 463894
rect 346584 463830 346636 463836
rect 346492 463140 346544 463146
rect 346492 463082 346544 463088
rect 345756 460080 345808 460086
rect 345756 460022 345808 460028
rect 345386 458552 345442 458561
rect 345386 458487 345442 458496
rect 343652 456766 343956 456794
rect 343824 453416 343876 453422
rect 343824 453358 343876 453364
rect 343180 453212 343232 453218
rect 343180 453154 343232 453160
rect 343192 449970 343220 453154
rect 342548 449942 342746 449970
rect 342824 449942 343114 449970
rect 343192 449942 343482 449970
rect 343836 449956 343864 453358
rect 343928 449970 343956 456766
rect 344560 454640 344612 454646
rect 344560 454582 344612 454588
rect 343928 449942 344218 449970
rect 344572 449956 344600 454582
rect 344926 450800 344982 450809
rect 344926 450735 344982 450744
rect 344940 449956 344968 450735
rect 345296 450152 345348 450158
rect 345296 450094 345348 450100
rect 345308 449956 345336 450094
rect 345400 449970 345428 458487
rect 345768 449970 345796 460022
rect 346504 449970 346532 463082
rect 346596 460934 346624 463830
rect 347780 461508 347832 461514
rect 347780 461450 347832 461456
rect 347792 460934 347820 461450
rect 346596 460906 346900 460934
rect 347792 460906 348740 460934
rect 346768 450356 346820 450362
rect 346768 450298 346820 450304
rect 345400 449942 345690 449970
rect 345768 449942 346058 449970
rect 346426 449942 346532 449970
rect 346780 449956 346808 450298
rect 346872 449970 346900 460906
rect 348330 459096 348386 459105
rect 348330 459031 348386 459040
rect 347964 458992 348016 458998
rect 347964 458934 348016 458940
rect 347504 454572 347556 454578
rect 347504 454514 347556 454520
rect 346872 449942 347162 449970
rect 347516 449956 347544 454514
rect 347872 453688 347924 453694
rect 347872 453630 347924 453636
rect 347884 449956 347912 453630
rect 347976 449970 348004 458934
rect 348056 456884 348108 456890
rect 348056 456826 348108 456832
rect 348068 453694 348096 456826
rect 348056 453688 348108 453694
rect 348056 453630 348108 453636
rect 348344 449970 348372 459031
rect 348712 449970 348740 460906
rect 349172 453218 349200 464063
rect 354678 463992 354734 464001
rect 354678 463927 354734 463936
rect 349252 463208 349304 463214
rect 349252 463150 349304 463156
rect 349160 453212 349212 453218
rect 349160 453154 349212 453160
rect 349264 449970 349292 463150
rect 351920 462528 351972 462534
rect 351920 462470 351972 462476
rect 351932 460934 351960 462470
rect 351932 460906 352788 460934
rect 350908 459944 350960 459950
rect 350908 459886 350960 459892
rect 349804 453212 349856 453218
rect 349804 453154 349856 453160
rect 349712 452192 349764 452198
rect 349712 452134 349764 452140
rect 347976 449942 348266 449970
rect 348344 449942 348634 449970
rect 348712 449942 349002 449970
rect 349264 449942 349370 449970
rect 349724 449956 349752 452134
rect 349816 449970 349844 453154
rect 350448 451104 350500 451110
rect 350448 451046 350500 451052
rect 349816 449942 350106 449970
rect 350460 449956 350488 451046
rect 350814 450664 350870 450673
rect 350814 450599 350870 450608
rect 350828 449956 350856 450599
rect 350920 449970 350948 459886
rect 352380 456068 352432 456074
rect 352380 456010 352432 456016
rect 352286 451888 352342 451897
rect 352286 451823 352342 451832
rect 351550 450256 351606 450265
rect 351550 450191 351606 450200
rect 351920 450220 351972 450226
rect 350920 449942 351210 449970
rect 351564 449956 351592 450191
rect 351920 450162 351972 450168
rect 351932 449956 351960 450162
rect 352300 449956 352328 451823
rect 352392 449970 352420 456010
rect 352760 449970 352788 460906
rect 353852 459060 353904 459066
rect 353852 459002 353904 459008
rect 353300 454504 353352 454510
rect 353300 454446 353352 454452
rect 353312 449970 353340 454446
rect 353758 450392 353814 450401
rect 353758 450327 353814 450336
rect 352392 449942 352682 449970
rect 352760 449942 353050 449970
rect 353312 449942 353418 449970
rect 353772 449956 353800 450327
rect 353864 449970 353892 459002
rect 354220 457632 354272 457638
rect 354220 457574 354272 457580
rect 354232 449970 354260 457574
rect 354692 456142 354720 463927
rect 358818 463856 358874 463865
rect 358818 463791 358874 463800
rect 354772 462528 354824 462534
rect 354772 462470 354824 462476
rect 354784 460934 354812 462470
rect 357440 461440 357492 461446
rect 357440 461382 357492 461388
rect 354784 460906 354996 460934
rect 354864 460624 354916 460630
rect 354864 460566 354916 460572
rect 354680 456136 354732 456142
rect 354680 456078 354732 456084
rect 353864 449942 354154 449970
rect 354232 449942 354522 449970
rect 354876 449956 354904 460566
rect 354968 449970 354996 460906
rect 356796 460080 356848 460086
rect 356796 460022 356848 460028
rect 356428 457700 356480 457706
rect 356428 457642 356480 457648
rect 355692 456136 355744 456142
rect 355692 456078 355744 456084
rect 355704 449970 355732 456078
rect 356060 453144 356112 453150
rect 356060 453086 356112 453092
rect 356072 449970 356100 453086
rect 356440 449970 356468 457642
rect 356808 449970 356836 460022
rect 357346 450936 357402 450945
rect 357346 450871 357402 450880
rect 357360 449970 357388 450871
rect 357452 450106 357480 461382
rect 357898 456920 357954 456929
rect 357898 456855 357954 456864
rect 357452 450078 357572 450106
rect 357544 449970 357572 450078
rect 357912 449970 357940 456855
rect 358268 455728 358320 455734
rect 358268 455670 358320 455676
rect 358280 449970 358308 455670
rect 358728 450560 358780 450566
rect 358728 450502 358780 450508
rect 358740 450265 358768 450502
rect 358726 450256 358782 450265
rect 358726 450191 358782 450200
rect 358832 449970 358860 463791
rect 361578 463720 361634 463729
rect 361578 463655 361634 463664
rect 360290 460048 360346 460057
rect 360290 459983 360346 459992
rect 359004 457768 359056 457774
rect 359004 457710 359056 457716
rect 359016 449970 359044 457710
rect 359372 457564 359424 457570
rect 359372 457506 359424 457512
rect 359384 449970 359412 457506
rect 360014 451480 360070 451489
rect 360014 451415 360070 451424
rect 354968 449942 355258 449970
rect 355704 449942 355994 449970
rect 356072 449942 356362 449970
rect 356440 449942 356730 449970
rect 356808 449942 357098 449970
rect 357360 449942 357466 449970
rect 357544 449942 357834 449970
rect 357912 449942 358202 449970
rect 358280 449942 358570 449970
rect 358832 449942 358938 449970
rect 359016 449942 359306 449970
rect 359384 449942 359674 449970
rect 360028 449956 360056 451415
rect 360198 450120 360254 450129
rect 360304 450106 360332 459983
rect 360842 455968 360898 455977
rect 360842 455903 360898 455912
rect 360304 450078 360516 450106
rect 360198 450055 360254 450064
rect 360212 449970 360240 450055
rect 360488 449970 360516 450078
rect 360856 449970 360884 455903
rect 361212 454504 361264 454510
rect 361212 454446 361264 454452
rect 361224 449970 361252 454446
rect 361592 449970 361620 463655
rect 364338 462360 364394 462369
rect 364338 462295 364394 462304
rect 362960 461372 363012 461378
rect 362960 461314 363012 461320
rect 361948 457836 362000 457842
rect 361948 457778 362000 457784
rect 361960 449970 361988 457778
rect 362972 450294 363000 461314
rect 364352 460934 364380 462295
rect 367112 460934 367140 465462
rect 370136 465452 370188 465458
rect 370136 465394 370188 465400
rect 368480 461304 368532 461310
rect 368480 461246 368532 461252
rect 368492 460934 368520 461246
rect 370148 460934 370176 465394
rect 372620 465384 372672 465390
rect 372620 465326 372672 465332
rect 371238 461408 371294 461417
rect 371238 461343 371294 461352
rect 371252 460934 371280 461343
rect 372632 460934 372660 465326
rect 375380 465316 375432 465322
rect 375380 465258 375432 465264
rect 364352 460906 364564 460934
rect 367112 460906 367508 460934
rect 368492 460906 369348 460934
rect 370148 460906 370452 460934
rect 371252 460906 371924 460934
rect 372632 460906 373396 460934
rect 363786 455832 363842 455841
rect 363786 455767 363842 455776
rect 363234 455560 363290 455569
rect 363234 455495 363290 455504
rect 363144 454572 363196 454578
rect 363144 454514 363196 454520
rect 362960 450288 363012 450294
rect 362960 450230 363012 450236
rect 362592 450220 362644 450226
rect 362592 450162 362644 450168
rect 360212 449942 360410 449970
rect 360488 449942 360778 449970
rect 360856 449942 361146 449970
rect 361224 449942 361514 449970
rect 361592 449942 361882 449970
rect 361960 449942 362250 449970
rect 362604 449956 362632 450162
rect 363156 449970 363184 454514
rect 362986 449942 363184 449970
rect 363248 449970 363276 455495
rect 363420 450288 363472 450294
rect 363420 450230 363472 450236
rect 363432 449970 363460 450230
rect 363800 449970 363828 455767
rect 364340 453144 364392 453150
rect 364340 453086 364392 453092
rect 364352 449970 364380 453086
rect 364536 449970 364564 460906
rect 366362 459912 366418 459921
rect 366362 459847 366418 459856
rect 364892 456816 364944 456822
rect 364892 456758 364944 456764
rect 364904 449970 364932 456758
rect 365994 456376 366050 456385
rect 365994 456311 366050 456320
rect 365904 450560 365956 450566
rect 365904 450502 365956 450508
rect 365536 450492 365588 450498
rect 365536 450434 365588 450440
rect 363248 449942 363354 449970
rect 363432 449942 363722 449970
rect 363800 449942 364090 449970
rect 364352 449942 364458 449970
rect 364536 449942 364826 449970
rect 364904 449942 365194 449970
rect 365548 449956 365576 450434
rect 365916 449956 365944 450502
rect 366008 449970 366036 456311
rect 366376 449970 366404 459847
rect 366730 458280 366786 458289
rect 366730 458215 366786 458224
rect 366744 449970 366772 458215
rect 367376 452328 367428 452334
rect 367376 452270 367428 452276
rect 366008 449942 366298 449970
rect 366376 449942 366666 449970
rect 366744 449942 367034 449970
rect 367388 449956 367416 452270
rect 367480 449970 367508 460906
rect 368938 459232 368994 459241
rect 368938 459167 368994 459176
rect 367836 456408 367888 456414
rect 367836 456350 367888 456356
rect 367848 449970 367876 456350
rect 368664 455660 368716 455666
rect 368664 455602 368716 455608
rect 368676 449970 368704 455602
rect 368848 450696 368900 450702
rect 368848 450638 368900 450644
rect 367480 449942 367770 449970
rect 367848 449942 368138 449970
rect 368506 449942 368704 449970
rect 368860 449956 368888 450638
rect 368952 449970 368980 459167
rect 369320 449970 369348 460906
rect 369952 458244 370004 458250
rect 369952 458186 370004 458192
rect 368952 449942 369242 449970
rect 369320 449942 369610 449970
rect 369964 449956 369992 458186
rect 370320 452668 370372 452674
rect 370320 452610 370372 452616
rect 370332 449956 370360 452610
rect 370424 449970 370452 460906
rect 370780 456612 370832 456618
rect 370780 456554 370832 456560
rect 370792 449970 370820 456554
rect 371516 455592 371568 455598
rect 371516 455534 371568 455540
rect 371240 453348 371292 453354
rect 371240 453290 371292 453296
rect 371252 452198 371280 453290
rect 371240 452192 371292 452198
rect 371240 452134 371292 452140
rect 371424 450288 371476 450294
rect 371424 450230 371476 450236
rect 370424 449942 370714 449970
rect 370792 449942 371082 449970
rect 371436 449956 371464 450230
rect 371528 449970 371556 455534
rect 371896 449970 371924 460906
rect 372250 459776 372306 459785
rect 372250 459711 372306 459720
rect 372264 449970 372292 459711
rect 372712 457632 372764 457638
rect 372712 457574 372764 457580
rect 372724 449970 372752 457574
rect 373264 451308 373316 451314
rect 373264 451250 373316 451256
rect 371528 449942 371818 449970
rect 371896 449942 372186 449970
rect 372264 449942 372554 449970
rect 372724 449942 372922 449970
rect 373276 449956 373304 451250
rect 373368 449970 373396 460906
rect 375288 456816 375340 456822
rect 375288 456758 375340 456764
rect 374092 456476 374144 456482
rect 374092 456418 374144 456424
rect 374104 449970 374132 456418
rect 374460 455796 374512 455802
rect 374460 455738 374512 455744
rect 373368 449942 373658 449970
rect 374026 449942 374132 449970
rect 374276 450016 374328 450022
rect 374472 449970 374500 455738
rect 375300 453354 375328 456758
rect 375392 456142 375420 465258
rect 380900 463820 380952 463826
rect 380900 463762 380952 463768
rect 378140 463344 378192 463350
rect 378140 463286 378192 463292
rect 375472 462596 375524 462602
rect 375472 462538 375524 462544
rect 375380 456136 375432 456142
rect 375380 456078 375432 456084
rect 375288 453348 375340 453354
rect 375288 453290 375340 453296
rect 375196 452328 375248 452334
rect 375196 452270 375248 452276
rect 375208 451382 375236 452270
rect 375196 451376 375248 451382
rect 375196 451318 375248 451324
rect 375104 450900 375156 450906
rect 375104 450842 375156 450848
rect 374328 449964 374394 449970
rect 374276 449958 374394 449964
rect 374288 449942 374394 449958
rect 374472 449942 374762 449970
rect 375116 449956 375144 450842
rect 375484 449956 375512 462538
rect 377034 461272 377090 461281
rect 377034 461207 377090 461216
rect 377048 460934 377076 461207
rect 377048 460906 377812 460934
rect 377036 456340 377088 456346
rect 377036 456282 377088 456288
rect 376300 456136 376352 456142
rect 376300 456078 376352 456084
rect 376392 456136 376444 456142
rect 376392 456078 376444 456084
rect 375932 454164 375984 454170
rect 375932 454106 375984 454112
rect 375838 451752 375894 451761
rect 375838 451687 375894 451696
rect 375852 449956 375880 451687
rect 375944 449970 375972 454106
rect 376312 449970 376340 456078
rect 376404 455802 376432 456078
rect 376392 455796 376444 455802
rect 376392 455738 376444 455744
rect 376760 455524 376812 455530
rect 376760 455466 376812 455472
rect 376772 449970 376800 455466
rect 377048 449970 377076 456282
rect 377404 455524 377456 455530
rect 377404 455466 377456 455472
rect 377416 449970 377444 455466
rect 377784 449970 377812 460906
rect 378152 449970 378180 463286
rect 380912 456794 380940 463762
rect 380990 461136 381046 461145
rect 380990 461071 381046 461080
rect 381004 460934 381032 461071
rect 383658 461000 383714 461009
rect 383658 460935 383714 460944
rect 381004 460906 381216 460934
rect 380912 456766 381124 456794
rect 379518 455560 379574 455569
rect 379518 455495 379574 455504
rect 378784 452192 378836 452198
rect 378784 452134 378836 452140
rect 378796 451858 378824 452134
rect 378784 451852 378836 451858
rect 378784 451794 378836 451800
rect 378782 450120 378838 450129
rect 378782 450055 378838 450064
rect 375944 449942 376234 449970
rect 376312 449942 376602 449970
rect 376772 449942 376970 449970
rect 377048 449942 377338 449970
rect 377416 449942 377706 449970
rect 377784 449942 378074 449970
rect 378152 449942 378442 449970
rect 378796 449956 378824 450055
rect 379532 449956 379560 455495
rect 379888 455456 379940 455462
rect 379888 455398 379940 455404
rect 379900 449956 379928 455398
rect 380254 452840 380310 452849
rect 380254 452775 380310 452784
rect 380268 449956 380296 452775
rect 380992 451852 381044 451858
rect 380992 451794 381044 451800
rect 380650 449954 380848 449970
rect 381004 449956 381032 451794
rect 381096 449970 381124 456766
rect 381188 451858 381216 460906
rect 382556 459672 382608 459678
rect 382556 459614 382608 459620
rect 381728 455456 381780 455462
rect 381728 455398 381780 455404
rect 381176 451852 381228 451858
rect 381176 451794 381228 451800
rect 380650 449948 380860 449954
rect 380650 449942 380808 449948
rect 279054 449919 279110 449928
rect 278504 449890 278556 449896
rect 381096 449942 381386 449970
rect 381740 449956 381768 455398
rect 382186 452976 382242 452985
rect 382186 452911 382242 452920
rect 382200 450634 382228 452911
rect 382188 450628 382240 450634
rect 382188 450570 382240 450576
rect 382568 449970 382596 459614
rect 383474 454064 383530 454073
rect 383474 453999 383530 454008
rect 383488 451897 383516 453999
rect 383566 452160 383622 452169
rect 383566 452095 383622 452104
rect 383474 451888 383530 451897
rect 383474 451823 383530 451832
rect 383476 450084 383528 450090
rect 383476 450026 383528 450032
rect 383488 449970 383516 450026
rect 382568 449942 382858 449970
rect 383226 449942 383516 449970
rect 383580 449956 383608 452095
rect 383672 449970 383700 460935
rect 385500 459740 385552 459746
rect 385500 459682 385552 459688
rect 384304 454096 384356 454102
rect 384304 454038 384356 454044
rect 383672 449942 383962 449970
rect 384316 449956 384344 454038
rect 385040 452328 385092 452334
rect 385040 452270 385092 452276
rect 384670 451888 384726 451897
rect 384670 451823 384726 451832
rect 384684 449956 384712 451823
rect 385052 449956 385080 452270
rect 385224 452192 385276 452198
rect 385224 452134 385276 452140
rect 380808 449890 380860 449896
rect 252586 449806 252876 449834
rect 355598 449848 355654 449857
rect 229742 449783 229798 449792
rect 382122 449818 382320 449834
rect 382122 449812 382332 449818
rect 382122 449806 382280 449812
rect 355598 449783 355654 449792
rect 382280 449754 382332 449760
rect 228088 449744 228140 449750
rect 382740 449744 382792 449750
rect 228140 449692 228298 449698
rect 228088 449686 228298 449692
rect 228100 449670 228298 449686
rect 379178 449682 379468 449698
rect 382490 449692 382740 449698
rect 382490 449686 382792 449692
rect 379178 449676 379480 449682
rect 379178 449670 379428 449676
rect 382490 449670 382780 449686
rect 379428 449618 379480 449624
rect 385236 449614 385264 452134
rect 385512 449970 385540 459682
rect 388904 456816 388956 456822
rect 388904 456758 388956 456764
rect 388536 454912 388588 454918
rect 388536 454854 388588 454860
rect 387708 452260 387760 452266
rect 387708 452202 387760 452208
rect 385512 449942 385802 449970
rect 386340 449806 386552 449834
rect 386142 449712 386198 449721
rect 386340 449698 386368 449806
rect 386524 449750 386552 449806
rect 387720 449750 387748 452202
rect 388442 450800 388498 450809
rect 388442 450735 388498 450744
rect 386420 449744 386472 449750
rect 386198 449670 386368 449698
rect 386418 449712 386420 449721
rect 386512 449744 386564 449750
rect 386472 449712 386474 449721
rect 386142 449647 386198 449656
rect 386512 449686 386564 449692
rect 387616 449744 387668 449750
rect 387616 449686 387668 449692
rect 387708 449744 387760 449750
rect 387708 449686 387760 449692
rect 386418 449647 386474 449656
rect 200856 449608 200908 449614
rect 193218 449576 193274 449585
rect 193218 449511 193274 449520
rect 193954 449576 194010 449585
rect 200856 449550 200908 449556
rect 201224 449608 201276 449614
rect 201224 449550 201276 449556
rect 307208 449608 307260 449614
rect 336740 449608 336792 449614
rect 307260 449556 307418 449562
rect 307208 449550 307418 449556
rect 385224 449608 385276 449614
rect 336792 449556 336858 449562
rect 336740 449550 336858 449556
rect 385684 449608 385736 449614
rect 385224 449550 385276 449556
rect 385434 449556 385684 449562
rect 387628 449585 387656 449686
rect 388076 449608 388128 449614
rect 385434 449550 385736 449556
rect 387614 449576 387670 449585
rect 307220 449534 307418 449550
rect 336752 449534 336858 449550
rect 385434 449534 385724 449550
rect 193954 449511 194010 449520
rect 388076 449550 388128 449556
rect 387614 449511 387670 449520
rect 194046 449304 194102 449313
rect 194046 449239 194102 449248
rect 191838 345128 191894 345137
rect 191838 345063 191894 345072
rect 190748 344986 191144 345014
rect 191116 147014 191144 344986
rect 388088 267734 388116 449550
rect 388088 267706 388300 267734
rect 388168 251864 388220 251870
rect 388168 251806 388220 251812
rect 388180 250730 388208 251806
rect 387918 250702 388208 250730
rect 308586 250472 308642 250481
rect 308586 250407 308642 250416
rect 191944 244934 191972 250036
rect 193232 250022 193338 250050
rect 194612 250022 194718 250050
rect 191932 244928 191984 244934
rect 191932 244870 191984 244876
rect 193232 233918 193260 250022
rect 193220 233912 193272 233918
rect 193220 233854 193272 233860
rect 191104 147008 191156 147014
rect 191104 146950 191156 146956
rect 190460 86284 190512 86290
rect 190460 86226 190512 86232
rect 190368 6860 190420 6866
rect 190368 6802 190420 6808
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 86226
rect 194612 39370 194640 250022
rect 196084 247110 196112 250036
rect 195244 247104 195296 247110
rect 195244 247046 195296 247052
rect 196072 247104 196124 247110
rect 196072 247046 196124 247052
rect 194600 39364 194652 39370
rect 194600 39306 194652 39312
rect 194416 4888 194468 4894
rect 194416 4830 194468 4836
rect 194428 480 194456 4830
rect 195256 4826 195284 247046
rect 197360 233912 197412 233918
rect 197360 233854 197412 233860
rect 197372 16574 197400 233854
rect 197464 42090 197492 250036
rect 198752 250022 198858 250050
rect 197452 42084 197504 42090
rect 197452 42026 197504 42032
rect 197372 16546 197952 16574
rect 195244 4820 195296 4826
rect 195244 4762 195296 4768
rect 197924 480 197952 16546
rect 198752 7614 198780 250022
rect 200224 247110 200252 250036
rect 201512 250022 201618 250050
rect 202892 250022 202998 250050
rect 204272 250022 204378 250050
rect 205652 250022 205758 250050
rect 207032 250022 207138 250050
rect 208412 250022 208518 250050
rect 209792 250022 209898 250050
rect 211172 250022 211278 250050
rect 199384 247104 199436 247110
rect 199384 247046 199436 247052
rect 200212 247104 200264 247110
rect 200212 247046 200264 247052
rect 199396 46238 199424 247046
rect 199384 46232 199436 46238
rect 199384 46174 199436 46180
rect 201512 16574 201540 250022
rect 201512 16546 201632 16574
rect 198740 7608 198792 7614
rect 198740 7550 198792 7556
rect 201500 7608 201552 7614
rect 201500 7550 201552 7556
rect 201512 480 201540 7550
rect 201604 3466 201632 16546
rect 202892 3534 202920 250022
rect 204272 3602 204300 250022
rect 205652 3670 205680 250022
rect 207032 3738 207060 250022
rect 208412 3806 208440 250022
rect 209792 3874 209820 250022
rect 211172 89010 211200 250022
rect 212644 245002 212672 250036
rect 213932 250022 214038 250050
rect 215312 250022 215418 250050
rect 216692 250022 216798 250050
rect 218072 250022 218178 250050
rect 219452 250022 219558 250050
rect 212632 244996 212684 245002
rect 212632 244938 212684 244944
rect 211160 89004 211212 89010
rect 211160 88946 211212 88952
rect 211160 24132 211212 24138
rect 211160 24074 211212 24080
rect 211172 16574 211200 24074
rect 211172 16546 211752 16574
rect 209780 3868 209832 3874
rect 209780 3810 209832 3816
rect 208400 3800 208452 3806
rect 208400 3742 208452 3748
rect 207020 3732 207072 3738
rect 207020 3674 207072 3680
rect 205640 3664 205692 3670
rect 205640 3606 205692 3612
rect 204260 3596 204312 3602
rect 204260 3538 204312 3544
rect 202880 3528 202932 3534
rect 202880 3470 202932 3476
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 201592 3460 201644 3466
rect 201592 3402 201644 3408
rect 205088 3460 205140 3466
rect 205088 3402 205140 3408
rect 205100 480 205128 3402
rect 208596 480 208624 3470
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213932 8974 213960 250022
rect 215312 228410 215340 250022
rect 215300 228404 215352 228410
rect 215300 228346 215352 228352
rect 216692 227050 216720 250022
rect 218072 240786 218100 250022
rect 218704 247716 218756 247722
rect 218704 247658 218756 247664
rect 218060 240780 218112 240786
rect 218060 240722 218112 240728
rect 216680 227044 216732 227050
rect 216680 226986 216732 226992
rect 213920 8968 213972 8974
rect 213920 8910 213972 8916
rect 215668 3596 215720 3602
rect 215668 3538 215720 3544
rect 215680 480 215708 3538
rect 218716 3466 218744 247658
rect 219452 225622 219480 250022
rect 220084 247852 220136 247858
rect 220084 247794 220136 247800
rect 219440 225616 219492 225622
rect 219440 225558 219492 225564
rect 219256 3664 219308 3670
rect 219256 3606 219308 3612
rect 218704 3460 218756 3466
rect 218704 3402 218756 3408
rect 219268 480 219296 3606
rect 220096 3534 220124 247794
rect 220924 242214 220952 250036
rect 222212 250022 222318 250050
rect 223592 250022 223698 250050
rect 224972 250022 225078 250050
rect 226352 250022 226458 250050
rect 220912 242208 220964 242214
rect 220912 242150 220964 242156
rect 222212 86290 222240 250022
rect 222844 247784 222896 247790
rect 222844 247726 222896 247732
rect 222200 86284 222252 86290
rect 222200 86226 222252 86232
rect 222856 3602 222884 247726
rect 223592 4894 223620 250022
rect 224224 247920 224276 247926
rect 224224 247862 224276 247868
rect 223580 4888 223632 4894
rect 223580 4830 223632 4836
rect 224236 3670 224264 247862
rect 224972 233918 225000 250022
rect 224960 233912 225012 233918
rect 224960 233854 225012 233860
rect 226352 7614 226380 250022
rect 227824 247722 227852 250036
rect 229204 247858 229232 250036
rect 230492 250022 230598 250050
rect 229192 247852 229244 247858
rect 229192 247794 229244 247800
rect 227812 247716 227864 247722
rect 227812 247658 227864 247664
rect 228364 247716 228416 247722
rect 228364 247658 228416 247664
rect 226340 7608 226392 7614
rect 226340 7550 226392 7556
rect 224224 3664 224276 3670
rect 224224 3606 224276 3612
rect 222844 3596 222896 3602
rect 222844 3538 222896 3544
rect 228376 3534 228404 247658
rect 230492 24138 230520 250022
rect 231964 247790 231992 250036
rect 233344 247926 233372 250036
rect 234632 250022 234738 250050
rect 233332 247920 233384 247926
rect 233332 247862 233384 247868
rect 231952 247784 232004 247790
rect 231952 247726 232004 247732
rect 234632 87378 234660 250022
rect 236104 247722 236132 250036
rect 237392 250022 237498 250050
rect 238772 250022 238878 250050
rect 236092 247716 236144 247722
rect 236092 247658 236144 247664
rect 233884 87372 233936 87378
rect 233884 87314 233936 87320
rect 234620 87372 234672 87378
rect 234620 87314 234672 87320
rect 230480 24132 230532 24138
rect 230480 24074 230532 24080
rect 220084 3528 220136 3534
rect 220084 3470 220136 3476
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 228364 3528 228416 3534
rect 228364 3470 228416 3476
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 222752 3460 222804 3466
rect 222752 3402 222804 3408
rect 222764 480 222792 3402
rect 226352 480 226380 3470
rect 229848 480 229876 3470
rect 233896 3466 233924 87314
rect 237392 3534 237420 250022
rect 237380 3528 237432 3534
rect 237380 3470 237432 3476
rect 233884 3460 233936 3466
rect 233884 3402 233936 3408
rect 238772 3262 238800 250022
rect 240244 247110 240272 250036
rect 241532 250022 241638 250050
rect 242912 250022 243018 250050
rect 244292 250022 244398 250050
rect 245672 250022 245778 250050
rect 247052 250022 247158 250050
rect 248432 250022 248538 250050
rect 249812 250022 249918 250050
rect 251192 250022 251298 250050
rect 252572 250022 252678 250050
rect 253952 250022 254058 250050
rect 255332 250022 255438 250050
rect 256712 250022 256818 250050
rect 258092 250022 258198 250050
rect 259472 250022 259578 250050
rect 260852 250022 260958 250050
rect 262232 250022 262338 250050
rect 263612 250022 263718 250050
rect 264992 250022 265098 250050
rect 266372 250022 266478 250050
rect 267752 250022 267858 250050
rect 269132 250022 269238 250050
rect 270512 250022 270618 250050
rect 239404 247104 239456 247110
rect 239404 247046 239456 247052
rect 240232 247104 240284 247110
rect 240232 247046 240284 247052
rect 233424 3256 233476 3262
rect 233424 3198 233476 3204
rect 238760 3256 238812 3262
rect 238760 3198 238812 3204
rect 233436 480 233464 3198
rect 239416 3058 239444 247046
rect 241532 3534 241560 250022
rect 242912 3534 242940 250022
rect 244292 3602 244320 250022
rect 244280 3596 244332 3602
rect 244280 3538 244332 3544
rect 245672 3534 245700 250022
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241520 3528 241572 3534
rect 241520 3470 241572 3476
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 245660 3528 245712 3534
rect 245660 3470 245712 3476
rect 237012 3052 237064 3058
rect 237012 2994 237064 3000
rect 239404 3052 239456 3058
rect 239404 2994 239456 3000
rect 237024 480 237052 2994
rect 240520 480 240548 3470
rect 244108 480 244136 3470
rect 247052 3466 247080 250022
rect 248432 4010 248460 250022
rect 248420 4004 248472 4010
rect 248420 3946 248472 3952
rect 249812 3942 249840 250022
rect 249800 3936 249852 3942
rect 249800 3878 249852 3884
rect 251192 3874 251220 250022
rect 251180 3868 251232 3874
rect 251180 3810 251232 3816
rect 252572 3806 252600 250022
rect 252560 3800 252612 3806
rect 252560 3742 252612 3748
rect 253952 3738 253980 250022
rect 253940 3732 253992 3738
rect 253940 3674 253992 3680
rect 255332 3670 255360 250022
rect 255320 3664 255372 3670
rect 255320 3606 255372 3612
rect 256712 3602 256740 250022
rect 247592 3596 247644 3602
rect 247592 3538 247644 3544
rect 256700 3596 256752 3602
rect 256700 3538 256752 3544
rect 247040 3460 247092 3466
rect 247040 3402 247092 3408
rect 247604 480 247632 3538
rect 258092 3534 258120 250022
rect 258264 4004 258316 4010
rect 258264 3946 258316 3952
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 258080 3528 258132 3534
rect 258080 3470 258132 3476
rect 251192 480 251220 3470
rect 254676 3460 254728 3466
rect 254676 3402 254728 3408
rect 254688 480 254716 3402
rect 258276 480 258304 3946
rect 259472 3466 259500 250022
rect 260852 175982 260880 250022
rect 260840 175976 260892 175982
rect 260840 175918 260892 175924
rect 262232 8974 262260 250022
rect 262220 8968 262272 8974
rect 262220 8910 262272 8916
rect 263612 7682 263640 250022
rect 264992 180130 265020 250022
rect 264980 180124 265032 180130
rect 264980 180066 265032 180072
rect 266372 10334 266400 250022
rect 267752 87650 267780 250022
rect 269132 89010 269160 250022
rect 269120 89004 269172 89010
rect 269120 88946 269172 88952
rect 267740 87644 267792 87650
rect 267740 87586 267792 87592
rect 270512 11762 270540 250022
rect 271984 247110 272012 250036
rect 273272 250022 273378 250050
rect 274652 250022 274758 250050
rect 276032 250022 276138 250050
rect 277412 250022 277518 250050
rect 278792 250022 278898 250050
rect 280172 250022 280278 250050
rect 281552 250022 281658 250050
rect 282932 250022 283038 250050
rect 284312 250022 284418 250050
rect 285692 250022 285798 250050
rect 287072 250022 287178 250050
rect 288452 250022 288558 250050
rect 271972 247104 272024 247110
rect 271972 247046 272024 247052
rect 273272 14482 273300 250022
rect 273904 247104 273956 247110
rect 273904 247046 273956 247052
rect 273916 206310 273944 247046
rect 273904 206304 273956 206310
rect 273904 206246 273956 206252
rect 273260 14476 273312 14482
rect 273260 14418 273312 14424
rect 270500 11756 270552 11762
rect 270500 11698 270552 11704
rect 266360 10328 266412 10334
rect 266360 10270 266412 10276
rect 263600 7676 263652 7682
rect 263600 7618 263652 7624
rect 274652 5370 274680 250022
rect 274640 5364 274692 5370
rect 274640 5306 274692 5312
rect 276032 5302 276060 250022
rect 277412 7614 277440 250022
rect 277400 7608 277452 7614
rect 277400 7550 277452 7556
rect 276020 5296 276072 5302
rect 276020 5238 276072 5244
rect 278792 5234 278820 250022
rect 278780 5228 278832 5234
rect 278780 5170 278832 5176
rect 280172 5166 280200 250022
rect 280160 5160 280212 5166
rect 280160 5102 280212 5108
rect 281552 5098 281580 250022
rect 281540 5092 281592 5098
rect 281540 5034 281592 5040
rect 282932 5030 282960 250022
rect 282920 5024 282972 5030
rect 282920 4966 282972 4972
rect 284312 4962 284340 250022
rect 284300 4956 284352 4962
rect 284300 4898 284352 4904
rect 285692 4894 285720 250022
rect 285680 4888 285732 4894
rect 285680 4830 285732 4836
rect 287072 4826 287100 250022
rect 287704 175976 287756 175982
rect 287704 175918 287756 175924
rect 287060 4820 287112 4826
rect 287060 4762 287112 4768
rect 261760 3936 261812 3942
rect 261760 3878 261812 3884
rect 259460 3460 259512 3466
rect 259460 3402 259512 3408
rect 261772 480 261800 3878
rect 265348 3868 265400 3874
rect 265348 3810 265400 3816
rect 265360 480 265388 3810
rect 268844 3800 268896 3806
rect 268844 3742 268896 3748
rect 268856 480 268884 3742
rect 272432 3732 272484 3738
rect 272432 3674 272484 3680
rect 272444 480 272472 3674
rect 276020 3664 276072 3670
rect 276020 3606 276072 3612
rect 276032 480 276060 3606
rect 279516 3596 279568 3602
rect 279516 3538 279568 3544
rect 279528 480 279556 3538
rect 287716 3534 287744 175918
rect 288452 6254 288480 250022
rect 289924 247110 289952 250036
rect 291212 250022 291318 250050
rect 292592 250022 292698 250050
rect 293972 250022 294078 250050
rect 295352 250022 295458 250050
rect 296732 250022 296838 250050
rect 298112 250022 298218 250050
rect 289912 247104 289964 247110
rect 289912 247046 289964 247052
rect 288440 6248 288492 6254
rect 288440 6190 288492 6196
rect 291212 6186 291240 250022
rect 291936 8968 291988 8974
rect 291936 8910 291988 8916
rect 291200 6180 291252 6186
rect 291200 6122 291252 6128
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 287704 3528 287756 3534
rect 287704 3470 287756 3476
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 283116 480 283144 3470
rect 286600 3460 286652 3466
rect 286600 3402 286652 3408
rect 286612 480 286640 3402
rect 290200 480 290228 3470
rect 291948 3058 291976 8910
rect 292592 6594 292620 250022
rect 292580 6588 292632 6594
rect 292580 6530 292632 6536
rect 293972 6526 294000 250022
rect 294052 7676 294104 7682
rect 294052 7618 294104 7624
rect 293960 6520 294012 6526
rect 293960 6462 294012 6468
rect 291936 3052 291988 3058
rect 291936 2994 291988 3000
rect 293684 3052 293736 3058
rect 293684 2994 293736 3000
rect 293696 480 293724 2994
rect 294064 2922 294092 7618
rect 295352 6458 295380 250022
rect 296732 175982 296760 250022
rect 296720 175976 296772 175982
rect 296720 175918 296772 175924
rect 295340 6452 295392 6458
rect 295340 6394 295392 6400
rect 298112 4010 298140 250022
rect 299584 247110 299612 250036
rect 300872 250022 300978 250050
rect 302252 250022 302358 250050
rect 303632 250022 303738 250050
rect 305012 250022 305118 250050
rect 298744 247104 298796 247110
rect 298744 247046 298796 247052
rect 299572 247104 299624 247110
rect 299572 247046 299624 247052
rect 298756 15910 298784 247046
rect 299480 180124 299532 180130
rect 299480 180066 299532 180072
rect 298744 15904 298796 15910
rect 298744 15846 298796 15852
rect 298100 4004 298152 4010
rect 298100 3946 298152 3952
rect 299492 3534 299520 180066
rect 300872 6390 300900 250022
rect 302252 180130 302280 250022
rect 302884 247104 302936 247110
rect 302884 247046 302936 247052
rect 302240 180124 302292 180130
rect 302240 180066 302292 180072
rect 302896 86290 302924 247046
rect 303632 227050 303660 250022
rect 303620 227044 303672 227050
rect 303620 226986 303672 226992
rect 302884 86284 302936 86290
rect 302884 86226 302936 86232
rect 303896 10328 303948 10334
rect 303896 10270 303948 10276
rect 300860 6384 300912 6390
rect 300860 6326 300912 6332
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 294052 2916 294104 2922
rect 294052 2858 294104 2864
rect 297272 2916 297324 2922
rect 297272 2858 297324 2864
rect 297284 480 297312 2858
rect 300780 480 300808 3470
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 10270
rect 305012 3942 305040 250022
rect 306484 247858 306512 250036
rect 306472 247852 306524 247858
rect 306472 247794 306524 247800
rect 307864 247790 307892 250036
rect 308600 249422 308628 250407
rect 387996 250050 388024 250702
rect 308588 249416 308640 249422
rect 308588 249358 308640 249364
rect 307852 247784 307904 247790
rect 307852 247726 307904 247732
rect 309244 247722 309272 250036
rect 310532 250022 310638 250050
rect 309232 247716 309284 247722
rect 309232 247658 309284 247664
rect 309784 89004 309836 89010
rect 309784 88946 309836 88952
rect 305644 87644 305696 87650
rect 305644 87586 305696 87592
rect 305000 3936 305052 3942
rect 305000 3878 305052 3884
rect 305656 3738 305684 87586
rect 305644 3732 305696 3738
rect 305644 3674 305696 3680
rect 307944 3732 307996 3738
rect 307944 3674 307996 3680
rect 307956 480 307984 3674
rect 309796 3534 309824 88946
rect 310532 17270 310560 250022
rect 311164 249416 311216 249422
rect 311164 249358 311216 249364
rect 311176 235278 311204 249358
rect 312004 247110 312032 250036
rect 313292 250022 313398 250050
rect 314672 250022 314778 250050
rect 316052 250022 316158 250050
rect 317432 250022 317538 250050
rect 318812 250022 318918 250050
rect 320192 250022 320298 250050
rect 321572 250022 321678 250050
rect 322952 250022 323058 250050
rect 324332 250022 324438 250050
rect 311992 247104 312044 247110
rect 311992 247046 312044 247052
rect 311164 235272 311216 235278
rect 311164 235214 311216 235220
rect 313292 21418 313320 250022
rect 313924 247104 313976 247110
rect 313924 247046 313976 247052
rect 313936 35222 313964 247046
rect 313924 35216 313976 35222
rect 313924 35158 313976 35164
rect 314672 22778 314700 250022
rect 316052 37942 316080 250022
rect 316040 37936 316092 37942
rect 316040 37878 316092 37884
rect 317432 28286 317460 250022
rect 317512 206304 317564 206310
rect 317512 206246 317564 206252
rect 317420 28280 317472 28286
rect 317420 28222 317472 28228
rect 314660 22772 314712 22778
rect 314660 22714 314712 22720
rect 313280 21412 313332 21418
rect 313280 21354 313332 21360
rect 310520 17264 310572 17270
rect 310520 17206 310572 17212
rect 317524 16574 317552 206246
rect 318812 25566 318840 250022
rect 320192 29646 320220 250022
rect 321572 31074 321600 250022
rect 321560 31068 321612 31074
rect 321560 31010 321612 31016
rect 320180 29640 320232 29646
rect 320180 29582 320232 29588
rect 318800 25560 318852 25566
rect 318800 25502 318852 25508
rect 322952 24138 322980 250022
rect 322940 24132 322992 24138
rect 322940 24074 322992 24080
rect 317524 16546 318104 16574
rect 314660 11756 314712 11762
rect 314660 11698 314712 11704
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 311452 480 311480 3470
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 11698
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 322112 14476 322164 14482
rect 322112 14418 322164 14424
rect 322124 480 322152 14418
rect 324332 3874 324360 250022
rect 325804 247110 325832 250036
rect 327092 250022 327198 250050
rect 328472 250022 328578 250050
rect 329852 250022 329958 250050
rect 331232 250022 331338 250050
rect 325792 247104 325844 247110
rect 325792 247046 325844 247052
rect 325608 5364 325660 5370
rect 325608 5306 325660 5312
rect 324320 3868 324372 3874
rect 324320 3810 324372 3816
rect 325620 480 325648 5306
rect 327092 3806 327120 250022
rect 327080 3800 327132 3806
rect 327080 3742 327132 3748
rect 328472 3738 328500 250022
rect 329104 247104 329156 247110
rect 329104 247046 329156 247052
rect 329116 26926 329144 247046
rect 329104 26920 329156 26926
rect 329104 26862 329156 26868
rect 329196 5296 329248 5302
rect 329196 5238 329248 5244
rect 328460 3732 328512 3738
rect 328460 3674 328512 3680
rect 329208 480 329236 5238
rect 329852 3670 329880 250022
rect 329840 3664 329892 3670
rect 329840 3606 329892 3612
rect 331232 3602 331260 250022
rect 332704 247110 332732 250036
rect 333992 250022 334098 250050
rect 335372 250022 335478 250050
rect 336752 250022 336858 250050
rect 338132 250022 338238 250050
rect 339512 250022 339618 250050
rect 340892 250022 340998 250050
rect 342272 250022 342378 250050
rect 343652 250022 343758 250050
rect 345032 250022 345138 250050
rect 346412 250022 346518 250050
rect 347792 250022 347898 250050
rect 349172 250022 349278 250050
rect 350552 250022 350658 250050
rect 351932 250022 352038 250050
rect 353312 250022 353418 250050
rect 354692 250022 354798 250050
rect 356072 250022 356178 250050
rect 357452 250022 357558 250050
rect 358832 250022 358938 250050
rect 360212 250022 360318 250050
rect 361592 250022 361698 250050
rect 362972 250022 363078 250050
rect 364352 250022 364458 250050
rect 332692 247104 332744 247110
rect 332692 247046 332744 247052
rect 332692 7608 332744 7614
rect 332692 7550 332744 7556
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 332704 480 332732 7550
rect 333992 3534 334020 250022
rect 335372 7614 335400 250022
rect 336004 247104 336056 247110
rect 336004 247046 336056 247052
rect 336016 32434 336044 247046
rect 336752 43450 336780 250022
rect 336740 43444 336792 43450
rect 336740 43386 336792 43392
rect 336004 32428 336056 32434
rect 336004 32370 336056 32376
rect 338132 8974 338160 250022
rect 339512 10334 339540 250022
rect 340144 235272 340196 235278
rect 340144 235214 340196 235220
rect 340156 221134 340184 235214
rect 340144 221128 340196 221134
rect 340144 221070 340196 221076
rect 340892 44878 340920 250022
rect 340880 44872 340932 44878
rect 340880 44814 340932 44820
rect 342272 11762 342300 250022
rect 343652 39370 343680 250022
rect 343640 39364 343692 39370
rect 343640 39306 343692 39312
rect 345032 14482 345060 250022
rect 345112 221128 345164 221134
rect 345112 221070 345164 221076
rect 345124 214606 345152 221070
rect 345112 214600 345164 214606
rect 345112 214542 345164 214548
rect 345020 14476 345072 14482
rect 345020 14418 345072 14424
rect 346412 13122 346440 250022
rect 347792 42090 347820 250022
rect 347780 42084 347832 42090
rect 347780 42026 347832 42032
rect 346400 13116 346452 13122
rect 346400 13058 346452 13064
rect 342260 11756 342312 11762
rect 342260 11698 342312 11704
rect 339500 10328 339552 10334
rect 339500 10270 339552 10276
rect 338120 8968 338172 8974
rect 338120 8910 338172 8916
rect 335360 7608 335412 7614
rect 335360 7550 335412 7556
rect 349172 5302 349200 250022
rect 349160 5296 349212 5302
rect 349160 5238 349212 5244
rect 350552 5234 350580 250022
rect 351932 40730 351960 250022
rect 351920 40724 351972 40730
rect 351920 40666 351972 40672
rect 336280 5228 336332 5234
rect 336280 5170 336332 5176
rect 350540 5228 350592 5234
rect 350540 5170 350592 5176
rect 333980 3528 334032 3534
rect 333980 3470 334032 3476
rect 336292 480 336320 5170
rect 353312 5166 353340 250022
rect 339868 5160 339920 5166
rect 339868 5102 339920 5108
rect 353300 5160 353352 5166
rect 353300 5102 353352 5108
rect 339880 480 339908 5102
rect 354692 5098 354720 250022
rect 343364 5092 343416 5098
rect 343364 5034 343416 5040
rect 354680 5092 354732 5098
rect 354680 5034 354732 5040
rect 343376 480 343404 5034
rect 356072 5030 356100 250022
rect 346952 5024 347004 5030
rect 346952 4966 347004 4972
rect 356060 5024 356112 5030
rect 356060 4966 356112 4972
rect 346964 480 346992 4966
rect 357452 4962 357480 250022
rect 350448 4956 350500 4962
rect 350448 4898 350500 4904
rect 357440 4956 357492 4962
rect 357440 4898 357492 4904
rect 350460 480 350488 4898
rect 358832 4894 358860 250022
rect 359464 214600 359516 214606
rect 359464 214542 359516 214548
rect 359476 207670 359504 214542
rect 359464 207664 359516 207670
rect 359464 207606 359516 207612
rect 354036 4888 354088 4894
rect 354036 4830 354088 4836
rect 358820 4888 358872 4894
rect 358820 4830 358872 4836
rect 354048 480 354076 4830
rect 360212 4826 360240 250022
rect 361592 36582 361620 250022
rect 361580 36576 361632 36582
rect 361580 36518 361632 36524
rect 362972 6322 363000 250022
rect 364352 33794 364380 250022
rect 365824 246430 365852 250036
rect 367112 250022 367218 250050
rect 368492 250022 368598 250050
rect 369872 250022 369978 250050
rect 371252 250022 371358 250050
rect 365812 246424 365864 246430
rect 365812 246366 365864 246372
rect 364340 33788 364392 33794
rect 364340 33730 364392 33736
rect 367112 15910 367140 250022
rect 368492 238134 368520 250022
rect 368480 238128 368532 238134
rect 368480 238070 368532 238076
rect 364616 15904 364668 15910
rect 364616 15846 364668 15852
rect 367100 15904 367152 15910
rect 367100 15846 367152 15852
rect 362960 6316 363012 6322
rect 362960 6258 363012 6264
rect 361120 6248 361172 6254
rect 361120 6190 361172 6196
rect 357532 4820 357584 4826
rect 357532 4762 357584 4768
rect 360200 4820 360252 4826
rect 360200 4762 360252 4768
rect 357544 480 357572 4762
rect 361132 480 361160 6190
rect 364628 480 364656 15846
rect 369872 6254 369900 250022
rect 369860 6248 369912 6254
rect 369860 6190 369912 6196
rect 371252 6186 371280 250022
rect 372724 246362 372752 250036
rect 374012 250022 374118 250050
rect 375392 250022 375498 250050
rect 376772 250022 376878 250050
rect 387918 250036 388024 250050
rect 372712 246356 372764 246362
rect 372712 246298 372764 246304
rect 371700 6588 371752 6594
rect 371700 6530 371752 6536
rect 368204 6180 368256 6186
rect 368204 6122 368256 6128
rect 371240 6180 371292 6186
rect 371240 6122 371292 6128
rect 368216 480 368244 6122
rect 371712 480 371740 6530
rect 374012 3466 374040 250022
rect 375392 233918 375420 250022
rect 376772 236706 376800 250022
rect 378244 249762 378272 250036
rect 378232 249756 378284 249762
rect 378232 249698 378284 249704
rect 378784 249756 378836 249762
rect 378784 249698 378836 249704
rect 376760 236700 376812 236706
rect 376760 236642 376812 236648
rect 378796 235958 378824 249698
rect 379624 248402 379652 250036
rect 379612 248396 379664 248402
rect 379612 248338 379664 248344
rect 381004 248130 381032 250036
rect 382384 248402 382412 250036
rect 382372 248396 382424 248402
rect 382372 248338 382424 248344
rect 383764 248198 383792 250036
rect 385144 248402 385172 250036
rect 387904 250022 388024 250036
rect 385132 248396 385184 248402
rect 385132 248338 385184 248344
rect 383752 248192 383804 248198
rect 383752 248134 383804 248140
rect 380992 248124 381044 248130
rect 380992 248066 381044 248072
rect 387904 245682 387932 250022
rect 387064 245676 387116 245682
rect 387064 245618 387116 245624
rect 387892 245676 387944 245682
rect 387892 245618 387944 245624
rect 387076 240786 387104 245618
rect 387064 240780 387116 240786
rect 387064 240722 387116 240728
rect 378784 235952 378836 235958
rect 378784 235894 378836 235900
rect 375380 233912 375432 233918
rect 375380 233854 375432 233860
rect 387076 230450 387104 240722
rect 388272 238754 388300 267706
rect 388088 238726 388300 238754
rect 387064 230444 387116 230450
rect 387064 230386 387116 230392
rect 374644 207664 374696 207670
rect 374644 207606 374696 207612
rect 374656 170338 374684 207606
rect 382280 175976 382332 175982
rect 382280 175918 382332 175924
rect 374644 170332 374696 170338
rect 374644 170274 374696 170280
rect 377220 170332 377272 170338
rect 377220 170274 377272 170280
rect 377232 168026 377260 170274
rect 377220 168020 377272 168026
rect 377220 167962 377272 167968
rect 379520 168020 379572 168026
rect 379520 167962 379572 167968
rect 379532 164898 379560 167962
rect 379520 164892 379572 164898
rect 379520 164834 379572 164840
rect 382292 16574 382320 175918
rect 388088 48278 388116 238726
rect 388456 147393 388484 450735
rect 388548 347585 388576 454854
rect 388812 452940 388864 452946
rect 388812 452882 388864 452888
rect 388720 451648 388772 451654
rect 388720 451590 388772 451596
rect 388626 450664 388682 450673
rect 388626 450599 388682 450608
rect 388534 347576 388590 347585
rect 388534 347511 388590 347520
rect 388442 147384 388498 147393
rect 388442 147319 388498 147328
rect 388640 146577 388668 450599
rect 388732 364334 388760 451590
rect 388824 383654 388852 452882
rect 388916 385014 388944 456758
rect 388996 449744 389048 449750
rect 388996 449686 389048 449692
rect 389008 449546 389036 449686
rect 388996 449540 389048 449546
rect 388996 449482 389048 449488
rect 388904 385008 388956 385014
rect 388904 384950 388956 384956
rect 388824 383626 388944 383654
rect 388916 378826 388944 383626
rect 388904 378820 388956 378826
rect 388904 378762 388956 378768
rect 388732 364306 388944 364334
rect 388916 349110 388944 364306
rect 388904 349104 388956 349110
rect 388904 349046 388956 349052
rect 389192 248130 389220 678943
rect 389270 455560 389326 455569
rect 389270 455495 389326 455504
rect 389180 248124 389232 248130
rect 389180 248066 389232 248072
rect 388626 146568 388682 146577
rect 388626 146503 388682 146512
rect 389180 86284 389232 86290
rect 389180 86226 389232 86232
rect 388076 48272 388128 48278
rect 388076 48214 388128 48220
rect 389192 16574 389220 86226
rect 389284 49609 389312 455495
rect 389916 454844 389968 454850
rect 389916 454786 389968 454792
rect 389364 454096 389416 454102
rect 389364 454038 389416 454044
rect 389376 248305 389404 454038
rect 389824 451036 389876 451042
rect 389824 450978 389876 450984
rect 389362 248296 389418 248305
rect 389362 248231 389418 248240
rect 389836 248130 389864 450978
rect 389928 347138 389956 454786
rect 390284 453552 390336 453558
rect 390284 453494 390336 453500
rect 390192 453484 390244 453490
rect 390192 453426 390244 453432
rect 390100 453008 390152 453014
rect 390100 452950 390152 452956
rect 390006 449576 390062 449585
rect 390006 449511 390062 449520
rect 390020 359417 390048 449511
rect 390112 380186 390140 452950
rect 390204 381546 390232 453426
rect 390296 382974 390324 453494
rect 390376 385008 390428 385014
rect 390376 384950 390428 384956
rect 390284 382968 390336 382974
rect 390284 382910 390336 382916
rect 390192 381540 390244 381546
rect 390192 381482 390244 381488
rect 390100 380180 390152 380186
rect 390100 380122 390152 380128
rect 390006 359408 390062 359417
rect 390006 359343 390062 359352
rect 390388 349858 390416 384950
rect 390376 349852 390428 349858
rect 390376 349794 390428 349800
rect 389916 347132 389968 347138
rect 389916 347074 389968 347080
rect 389916 258120 389968 258126
rect 389916 258062 389968 258068
rect 389928 249762 389956 258062
rect 389916 249756 389968 249762
rect 389916 249698 389968 249704
rect 390572 248266 390600 681935
rect 390664 248402 390692 682479
rect 390742 682136 390798 682145
rect 390742 682071 390798 682080
rect 390652 248396 390704 248402
rect 390652 248338 390704 248344
rect 390560 248260 390612 248266
rect 390560 248202 390612 248208
rect 390756 248198 390784 682071
rect 396736 501634 396764 699654
rect 416778 536888 416834 536897
rect 406292 536852 406344 536858
rect 416778 536823 416780 536832
rect 406292 536794 406344 536800
rect 416832 536823 416834 536832
rect 416780 536794 416832 536800
rect 396724 501628 396776 501634
rect 396724 501570 396776 501576
rect 395344 464568 395396 464574
rect 395344 464510 395396 464516
rect 394056 464500 394108 464506
rect 394056 464442 394108 464448
rect 392952 455728 393004 455734
rect 392952 455670 393004 455676
rect 391296 454436 391348 454442
rect 391296 454378 391348 454384
rect 391204 454300 391256 454306
rect 391204 454242 391256 454248
rect 391216 347002 391244 454242
rect 391308 347546 391336 454378
rect 391388 454368 391440 454374
rect 391388 454310 391440 454316
rect 391400 347614 391428 454310
rect 392768 454164 392820 454170
rect 392768 454106 392820 454112
rect 392674 453384 392730 453393
rect 392674 453319 392730 453328
rect 392582 450392 392638 450401
rect 392582 450327 392638 450336
rect 391388 347608 391440 347614
rect 391388 347550 391440 347556
rect 391296 347540 391348 347546
rect 391296 347482 391348 347488
rect 391204 346996 391256 347002
rect 391204 346938 391256 346944
rect 390744 248192 390796 248198
rect 390744 248134 390796 248140
rect 389824 248124 389876 248130
rect 389824 248066 389876 248072
rect 392596 147529 392624 450327
rect 392688 259418 392716 453319
rect 392780 346322 392808 454106
rect 392860 452668 392912 452674
rect 392860 452610 392912 452616
rect 392768 346316 392820 346322
rect 392768 346258 392820 346264
rect 392872 346254 392900 452610
rect 392964 348498 392992 455670
rect 393962 453520 394018 453529
rect 393962 453455 394018 453464
rect 393136 453144 393188 453150
rect 393136 453086 393188 453092
rect 393044 451376 393096 451382
rect 393044 451318 393096 451324
rect 392952 348492 393004 348498
rect 392952 348434 393004 348440
rect 393056 348430 393084 451318
rect 393148 349178 393176 453086
rect 393136 349172 393188 349178
rect 393136 349114 393188 349120
rect 393044 348424 393096 348430
rect 393044 348366 393096 348372
rect 392860 346248 392912 346254
rect 392860 346190 392912 346196
rect 392676 259412 392728 259418
rect 392676 259354 392728 259360
rect 392582 147520 392638 147529
rect 392582 147455 392638 147464
rect 393976 59362 394004 453455
rect 394068 346050 394096 464442
rect 394332 455048 394384 455054
rect 394332 454990 394384 454996
rect 394148 454708 394200 454714
rect 394148 454650 394200 454656
rect 394056 346044 394108 346050
rect 394056 345986 394108 345992
rect 394160 345030 394188 454650
rect 394240 454232 394292 454238
rect 394240 454174 394292 454180
rect 394252 346186 394280 454174
rect 394240 346180 394292 346186
rect 394240 346122 394292 346128
rect 394344 345370 394372 454990
rect 394424 452328 394476 452334
rect 394424 452270 394476 452276
rect 394436 346390 394464 452270
rect 394516 451784 394568 451790
rect 394516 451726 394568 451732
rect 394424 346384 394476 346390
rect 394424 346326 394476 346332
rect 394528 345846 394556 451726
rect 394608 450764 394660 450770
rect 394608 450706 394660 450712
rect 394620 347682 394648 450706
rect 394608 347676 394660 347682
rect 394608 347618 394660 347624
rect 394516 345840 394568 345846
rect 394516 345782 394568 345788
rect 394332 345364 394384 345370
rect 394332 345306 394384 345312
rect 394148 345024 394200 345030
rect 394148 344966 394200 344972
rect 393964 59356 394016 59362
rect 393964 59298 394016 59304
rect 389270 49600 389326 49609
rect 389270 49535 389326 49544
rect 395356 46850 395384 464510
rect 406200 464296 406252 464302
rect 406200 464238 406252 464244
rect 395436 462868 395488 462874
rect 395436 462810 395488 462816
rect 395344 46844 395396 46850
rect 395344 46786 395396 46792
rect 395448 46714 395476 462810
rect 405004 462732 405056 462738
rect 405004 462674 405056 462680
rect 403624 462460 403676 462466
rect 403624 462402 403676 462408
rect 395528 461780 395580 461786
rect 395528 461722 395580 461728
rect 395540 46782 395568 461722
rect 400772 461576 400824 461582
rect 400772 461518 400824 461524
rect 396724 460012 396776 460018
rect 396724 459954 396776 459960
rect 395620 456068 395672 456074
rect 395620 456010 395672 456016
rect 395632 348634 395660 456010
rect 395804 453280 395856 453286
rect 395804 453222 395856 453228
rect 395712 450356 395764 450362
rect 395712 450298 395764 450304
rect 395620 348628 395672 348634
rect 395620 348570 395672 348576
rect 395724 347177 395752 450298
rect 395816 349314 395844 453222
rect 395896 453212 395948 453218
rect 395896 453154 395948 453160
rect 395908 349382 395936 453154
rect 395896 349376 395948 349382
rect 395896 349318 395948 349324
rect 395804 349308 395856 349314
rect 395804 349250 395856 349256
rect 395710 347168 395766 347177
rect 395710 347103 395766 347112
rect 396736 345710 396764 459954
rect 398104 456136 398156 456142
rect 398104 456078 398156 456084
rect 396816 454776 396868 454782
rect 396816 454718 396868 454724
rect 396828 345778 396856 454718
rect 397184 452124 397236 452130
rect 397184 452066 397236 452072
rect 397092 452056 397144 452062
rect 397092 451998 397144 452004
rect 396908 451988 396960 451994
rect 396908 451930 396960 451936
rect 396920 345982 396948 451930
rect 397000 451920 397052 451926
rect 397000 451862 397052 451868
rect 396908 345976 396960 345982
rect 396908 345918 396960 345924
rect 396816 345772 396868 345778
rect 396816 345714 396868 345720
rect 396724 345704 396776 345710
rect 396724 345646 396776 345652
rect 397012 345506 397040 451862
rect 397104 345642 397132 451998
rect 397196 345914 397224 452066
rect 397184 345908 397236 345914
rect 397184 345850 397236 345856
rect 397092 345636 397144 345642
rect 397092 345578 397144 345584
rect 397000 345500 397052 345506
rect 397000 345442 397052 345448
rect 398116 247217 398144 456078
rect 398196 455592 398248 455598
rect 398196 455534 398248 455540
rect 398208 249150 398236 455534
rect 398288 455524 398340 455530
rect 398288 455466 398340 455472
rect 398196 249144 398248 249150
rect 398196 249086 398248 249092
rect 398300 249082 398328 455466
rect 398656 453076 398708 453082
rect 398656 453018 398708 453024
rect 398378 452160 398434 452169
rect 398378 452095 398434 452104
rect 398288 249076 398340 249082
rect 398288 249018 398340 249024
rect 398102 247208 398158 247217
rect 398102 247143 398158 247152
rect 398392 247042 398420 452095
rect 398564 450696 398616 450702
rect 398564 450638 398616 450644
rect 398472 449948 398524 449954
rect 398472 449890 398524 449896
rect 398380 247036 398432 247042
rect 398380 246978 398432 246984
rect 398484 245614 398512 449890
rect 398576 246974 398604 450638
rect 398668 349450 398696 453018
rect 399484 449608 399536 449614
rect 399484 449550 399536 449556
rect 399496 349926 399524 449550
rect 399484 349920 399536 349926
rect 399484 349862 399536 349868
rect 400784 349518 400812 461518
rect 402520 460148 402572 460154
rect 402520 460090 402572 460096
rect 400956 460080 401008 460086
rect 400956 460022 401008 460028
rect 400864 459128 400916 459134
rect 400864 459070 400916 459076
rect 400772 349512 400824 349518
rect 400772 349454 400824 349460
rect 398656 349444 398708 349450
rect 398656 349386 398708 349392
rect 400876 248198 400904 459070
rect 400968 249354 400996 460022
rect 401048 459944 401100 459950
rect 401048 459886 401100 459892
rect 401060 249490 401088 459886
rect 402244 459876 402296 459882
rect 402244 459818 402296 459824
rect 401140 459060 401192 459066
rect 401140 459002 401192 459008
rect 401048 249484 401100 249490
rect 401048 249426 401100 249432
rect 401152 249422 401180 459002
rect 401232 458992 401284 458998
rect 401232 458934 401284 458940
rect 401244 249558 401272 458934
rect 401324 454572 401376 454578
rect 401324 454514 401376 454520
rect 401232 249552 401284 249558
rect 401232 249494 401284 249500
rect 401140 249416 401192 249422
rect 401140 249358 401192 249364
rect 400956 249348 401008 249354
rect 400956 249290 401008 249296
rect 401336 249218 401364 454514
rect 401506 451480 401562 451489
rect 401506 451415 401562 451424
rect 401416 450560 401468 450566
rect 401416 450502 401468 450508
rect 401324 249212 401376 249218
rect 401324 249154 401376 249160
rect 400864 248192 400916 248198
rect 400864 248134 400916 248140
rect 398564 246968 398616 246974
rect 398564 246910 398616 246916
rect 401428 246906 401456 450502
rect 401520 249286 401548 451415
rect 401508 249280 401560 249286
rect 401508 249222 401560 249228
rect 402256 248334 402284 459818
rect 402428 458924 402480 458930
rect 402428 458866 402480 458872
rect 402336 458788 402388 458794
rect 402336 458730 402388 458736
rect 402244 248328 402296 248334
rect 402244 248270 402296 248276
rect 402348 248266 402376 458730
rect 402336 248260 402388 248266
rect 402336 248202 402388 248208
rect 402440 248033 402468 458866
rect 402532 249665 402560 460090
rect 402612 458720 402664 458726
rect 402612 458662 402664 458668
rect 402518 249656 402574 249665
rect 402518 249591 402574 249600
rect 402426 248024 402482 248033
rect 402426 247959 402482 247968
rect 402624 247761 402652 458662
rect 403532 450424 403584 450430
rect 403532 450366 403584 450372
rect 403544 249762 403572 450366
rect 403532 249756 403584 249762
rect 403532 249698 403584 249704
rect 402610 247752 402666 247761
rect 402610 247687 402666 247696
rect 401416 246900 401468 246906
rect 401416 246842 401468 246848
rect 398472 245608 398524 245614
rect 398472 245550 398524 245556
rect 398840 227044 398892 227050
rect 398840 226986 398892 226992
rect 396080 180124 396132 180130
rect 396080 180066 396132 180072
rect 395528 46776 395580 46782
rect 395528 46718 395580 46724
rect 395436 46708 395488 46714
rect 395436 46650 395488 46656
rect 382292 16546 382412 16574
rect 389192 16546 389496 16574
rect 375288 6520 375340 6526
rect 375288 6462 375340 6468
rect 374000 3460 374052 3466
rect 374000 3402 374052 3408
rect 375300 480 375328 6462
rect 378876 6452 378928 6458
rect 378876 6394 378928 6400
rect 378888 480 378916 6394
rect 382384 480 382412 16546
rect 385960 4004 386012 4010
rect 385960 3946 386012 3952
rect 385972 480 386000 3946
rect 389468 480 389496 16546
rect 393044 6384 393096 6390
rect 393044 6326 393096 6332
rect 393056 480 393084 6326
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 180066
rect 398852 3398 398880 226986
rect 400864 164892 400916 164898
rect 400864 164834 400916 164840
rect 400876 158030 400904 164834
rect 400864 158024 400916 158030
rect 400864 157966 400916 157972
rect 403636 46646 403664 462402
rect 403992 458584 404044 458590
rect 403992 458526 404044 458532
rect 403900 458448 403952 458454
rect 403900 458390 403952 458396
rect 403806 456104 403862 456113
rect 403806 456039 403862 456048
rect 403716 456000 403768 456006
rect 403716 455942 403768 455948
rect 403728 149054 403756 455942
rect 403716 149048 403768 149054
rect 403716 148990 403768 148996
rect 403820 148986 403848 456039
rect 403912 245478 403940 458390
rect 404004 248169 404032 458526
rect 404084 458380 404136 458386
rect 404084 458322 404136 458328
rect 404096 249626 404124 458322
rect 404176 455932 404228 455938
rect 404176 455874 404228 455880
rect 404188 249694 404216 455874
rect 404268 450152 404320 450158
rect 404268 450094 404320 450100
rect 404176 249688 404228 249694
rect 404176 249630 404228 249636
rect 404084 249620 404136 249626
rect 404084 249562 404136 249568
rect 403990 248160 404046 248169
rect 403990 248095 404046 248104
rect 404280 245546 404308 450094
rect 404268 245540 404320 245546
rect 404268 245482 404320 245488
rect 403900 245472 403952 245478
rect 403900 245414 403952 245420
rect 403808 148980 403860 148986
rect 403808 148922 403860 148928
rect 405016 47977 405044 462674
rect 405372 460488 405424 460494
rect 405372 460430 405424 460436
rect 405280 460352 405332 460358
rect 405280 460294 405332 460300
rect 405094 458960 405150 458969
rect 405094 458895 405150 458904
rect 405108 48210 405136 458895
rect 405186 452976 405242 452985
rect 405186 452911 405242 452920
rect 405096 48204 405148 48210
rect 405096 48146 405148 48152
rect 405002 47968 405058 47977
rect 405002 47903 405058 47912
rect 405200 47841 405228 452911
rect 405292 247897 405320 460294
rect 405384 248946 405412 460430
rect 405464 458652 405516 458658
rect 405464 458594 405516 458600
rect 405476 249801 405504 458594
rect 406212 347449 406240 464238
rect 406198 347440 406254 347449
rect 406198 347375 406254 347384
rect 406304 251870 406332 536794
rect 416778 535936 416834 535945
rect 416778 535871 416834 535880
rect 416792 535498 416820 535871
rect 416780 535492 416832 535498
rect 416780 535434 416832 535440
rect 417054 533760 417110 533769
rect 417054 533695 417110 533704
rect 416044 532840 416096 532846
rect 416044 532782 416096 532788
rect 414664 530052 414716 530058
rect 414664 529994 414716 530000
rect 407856 463208 407908 463214
rect 407856 463150 407908 463156
rect 407764 462936 407816 462942
rect 407764 462878 407816 462884
rect 406842 457600 406898 457609
rect 406842 457535 406898 457544
rect 406658 457464 406714 457473
rect 406658 457399 406714 457408
rect 406474 457192 406530 457201
rect 406474 457127 406530 457136
rect 406382 454064 406438 454073
rect 406382 453999 406438 454008
rect 406292 251864 406344 251870
rect 406292 251806 406344 251812
rect 405462 249792 405518 249801
rect 405462 249727 405518 249736
rect 405372 248940 405424 248946
rect 405372 248882 405424 248888
rect 405278 247888 405334 247897
rect 405278 247823 405334 247832
rect 406396 49502 406424 453999
rect 406488 147626 406516 457127
rect 406568 457088 406620 457094
rect 406568 457030 406620 457036
rect 406580 148306 406608 457030
rect 406568 148300 406620 148306
rect 406568 148242 406620 148248
rect 406476 147620 406528 147626
rect 406476 147562 406528 147568
rect 406672 147558 406700 457399
rect 406750 455696 406806 455705
rect 406750 455631 406806 455640
rect 406764 148238 406792 455631
rect 406856 149297 406884 457535
rect 406934 452840 406990 452849
rect 406934 452775 406990 452784
rect 406842 149288 406898 149297
rect 406842 149223 406898 149232
rect 406948 148510 406976 452775
rect 407028 450084 407080 450090
rect 407028 450026 407080 450032
rect 406936 148504 406988 148510
rect 406936 148446 406988 148452
rect 407040 148442 407068 450026
rect 407120 247852 407172 247858
rect 407120 247794 407172 247800
rect 407028 148436 407080 148442
rect 407028 148378 407080 148384
rect 406752 148232 406804 148238
rect 406752 148174 406804 148180
rect 406660 147552 406712 147558
rect 406660 147494 406712 147500
rect 406384 49496 406436 49502
rect 406384 49438 406436 49444
rect 405186 47832 405242 47841
rect 405186 47767 405242 47776
rect 403624 46640 403676 46646
rect 403624 46582 403676 46588
rect 407132 16574 407160 247794
rect 407776 49473 407804 462878
rect 407868 49706 407896 463150
rect 410616 463140 410668 463146
rect 410616 463082 410668 463088
rect 408040 462800 408092 462806
rect 408040 462742 408092 462748
rect 407948 462664 408000 462670
rect 407948 462606 408000 462612
rect 407856 49700 407908 49706
rect 407856 49642 407908 49648
rect 407762 49464 407818 49473
rect 407762 49399 407818 49408
rect 407960 48890 407988 462606
rect 408052 49774 408080 462742
rect 410522 462496 410578 462505
rect 410522 462431 410578 462440
rect 408314 458824 408370 458833
rect 408314 458759 408370 458768
rect 408130 458416 408186 458425
rect 408130 458351 408186 458360
rect 408040 49768 408092 49774
rect 408040 49710 408092 49716
rect 408144 49337 408172 458351
rect 408222 453112 408278 453121
rect 408222 453047 408278 453056
rect 408236 349586 408264 453047
rect 408224 349580 408276 349586
rect 408224 349522 408276 349528
rect 408328 49842 408356 458759
rect 409142 457328 409198 457337
rect 409142 457263 409198 457272
rect 409156 147490 409184 457263
rect 409328 456340 409380 456346
rect 409328 456282 409380 456288
rect 409236 455660 409288 455666
rect 409236 455602 409288 455608
rect 409248 148714 409276 455602
rect 409236 148708 409288 148714
rect 409236 148650 409288 148656
rect 409340 148578 409368 456282
rect 409696 450968 409748 450974
rect 409696 450910 409748 450916
rect 409512 450492 409564 450498
rect 409512 450434 409564 450440
rect 409420 450288 409472 450294
rect 409420 450230 409472 450236
rect 409432 148646 409460 450230
rect 409524 148782 409552 450434
rect 409604 450016 409656 450022
rect 409604 449958 409656 449964
rect 409616 149122 409644 449958
rect 409708 347478 409736 450910
rect 409696 347472 409748 347478
rect 409696 347414 409748 347420
rect 409880 247784 409932 247790
rect 409880 247726 409932 247732
rect 409604 149116 409656 149122
rect 409604 149058 409656 149064
rect 409512 148776 409564 148782
rect 409512 148718 409564 148724
rect 409420 148640 409472 148646
rect 409420 148582 409472 148588
rect 409328 148572 409380 148578
rect 409328 148514 409380 148520
rect 409144 147484 409196 147490
rect 409144 147426 409196 147432
rect 408316 49836 408368 49842
rect 408316 49778 408368 49784
rect 408130 49328 408186 49337
rect 408130 49263 408186 49272
rect 407948 48884 408000 48890
rect 407948 48826 408000 48832
rect 409892 16574 409920 247726
rect 410536 48074 410564 462431
rect 410628 48958 410656 463082
rect 410708 463072 410760 463078
rect 410708 463014 410760 463020
rect 410720 49609 410748 463014
rect 413282 462632 413338 462641
rect 413282 462567 413338 462576
rect 410800 462528 410852 462534
rect 410800 462470 410852 462476
rect 410706 49600 410762 49609
rect 410812 49570 410840 462470
rect 411812 460420 411864 460426
rect 411812 460362 411864 460368
rect 410890 455968 410946 455977
rect 410890 455903 410946 455912
rect 410706 49535 410762 49544
rect 410800 49564 410852 49570
rect 410800 49506 410852 49512
rect 410904 49434 410932 455903
rect 410982 453248 411038 453257
rect 410982 453183 411038 453192
rect 410996 349217 411024 453183
rect 411076 449540 411128 449546
rect 411076 449482 411128 449488
rect 410982 349208 411038 349217
rect 410982 349143 411038 349152
rect 411088 348702 411116 449482
rect 411076 348696 411128 348702
rect 411076 348638 411128 348644
rect 411824 347342 411852 460362
rect 412364 457700 412416 457706
rect 412364 457642 412416 457648
rect 411996 457564 412048 457570
rect 411996 457506 412048 457512
rect 411902 450120 411958 450129
rect 411902 450055 411958 450064
rect 411812 347336 411864 347342
rect 411812 347278 411864 347284
rect 410984 158024 411036 158030
rect 410984 157966 411036 157972
rect 410996 148374 411024 157966
rect 410984 148368 411036 148374
rect 410984 148310 411036 148316
rect 410892 49428 410944 49434
rect 410892 49370 410944 49376
rect 411916 49094 411944 450055
rect 412008 148918 412036 457506
rect 412272 457360 412324 457366
rect 412272 457302 412324 457308
rect 412088 456952 412140 456958
rect 412088 456894 412140 456900
rect 412100 149326 412128 456894
rect 412180 456884 412232 456890
rect 412180 456826 412232 456832
rect 412088 149320 412140 149326
rect 412088 149262 412140 149268
rect 412192 149258 412220 456826
rect 412284 149462 412312 457302
rect 412272 149456 412324 149462
rect 412272 149398 412324 149404
rect 412180 149252 412232 149258
rect 412180 149194 412232 149200
rect 412376 149190 412404 457642
rect 412456 457428 412508 457434
rect 412456 457370 412508 457376
rect 412468 149394 412496 457370
rect 412548 450220 412600 450226
rect 412548 450162 412600 450168
rect 412456 149388 412508 149394
rect 412456 149330 412508 149336
rect 412364 149184 412416 149190
rect 412364 149126 412416 149132
rect 411996 148912 412048 148918
rect 411996 148854 412048 148860
rect 412560 148850 412588 450162
rect 412548 148844 412600 148850
rect 412548 148786 412600 148792
rect 411904 49088 411956 49094
rect 411904 49030 411956 49036
rect 410616 48952 410668 48958
rect 410616 48894 410668 48900
rect 413296 48142 413324 462567
rect 414676 461718 414704 529994
rect 416056 464438 416084 532782
rect 417068 532778 417096 533695
rect 418068 532840 418120 532846
rect 418066 532808 418068 532817
rect 418120 532808 418122 532817
rect 417056 532772 417108 532778
rect 418066 532743 418122 532752
rect 417056 532714 417108 532720
rect 417698 531040 417754 531049
rect 417698 530975 417754 530984
rect 417424 530052 417476 530058
rect 417424 529994 417476 530000
rect 417436 529961 417464 529994
rect 417712 529990 417740 530975
rect 417700 529984 417752 529990
rect 417422 529952 417478 529961
rect 417700 529926 417752 529932
rect 417422 529887 417478 529896
rect 417698 528184 417754 528193
rect 417698 528119 417754 528128
rect 417712 527202 417740 528119
rect 417700 527196 417752 527202
rect 417700 527138 417752 527144
rect 417606 509960 417662 509969
rect 417606 509895 417662 509904
rect 417620 509318 417648 509895
rect 417608 509312 417660 509318
rect 417608 509254 417660 509260
rect 418066 508328 418122 508337
rect 418066 508263 418122 508272
rect 416778 508056 416834 508065
rect 416778 507991 416834 508000
rect 416792 507890 416820 507991
rect 416780 507884 416832 507890
rect 416780 507826 416832 507832
rect 416044 464432 416096 464438
rect 416044 464374 416096 464380
rect 416044 462392 416096 462398
rect 416044 462334 416096 462340
rect 414664 461712 414716 461718
rect 414664 461654 414716 461660
rect 415308 458516 415360 458522
rect 415308 458458 415360 458464
rect 413466 458280 413522 458289
rect 413376 458244 413428 458250
rect 413466 458215 413522 458224
rect 413376 458186 413428 458192
rect 413388 49162 413416 458186
rect 413480 49298 413508 458215
rect 414664 457292 414716 457298
rect 414664 457234 414716 457240
rect 413558 456920 413614 456929
rect 413558 456855 413614 456864
rect 413572 49638 413600 456855
rect 414572 456544 414624 456550
rect 414572 456486 414624 456492
rect 413650 455832 413706 455841
rect 413650 455767 413706 455776
rect 413560 49632 413612 49638
rect 413560 49574 413612 49580
rect 413664 49366 413692 455767
rect 413836 451716 413888 451722
rect 413836 451658 413888 451664
rect 413744 451580 413796 451586
rect 413744 451522 413796 451528
rect 413756 346118 413784 451522
rect 413848 347274 413876 451658
rect 413928 449744 413980 449750
rect 413928 449686 413980 449692
rect 413940 348566 413968 449686
rect 414584 349042 414612 456486
rect 414572 349036 414624 349042
rect 414572 348978 414624 348984
rect 413928 348560 413980 348566
rect 413928 348502 413980 348508
rect 413836 347268 413888 347274
rect 413836 347210 413888 347216
rect 413744 346112 413796 346118
rect 413744 346054 413796 346060
rect 414572 345976 414624 345982
rect 414572 345918 414624 345924
rect 414480 345704 414532 345710
rect 414480 345646 414532 345652
rect 414020 247716 414072 247722
rect 414020 247658 414072 247664
rect 413652 49360 413704 49366
rect 413652 49302 413704 49308
rect 413468 49292 413520 49298
rect 413468 49234 413520 49240
rect 413376 49156 413428 49162
rect 413376 49098 413428 49104
rect 413284 48136 413336 48142
rect 413284 48078 413336 48084
rect 410524 48068 410576 48074
rect 410524 48010 410576 48016
rect 414032 16574 414060 247658
rect 414492 247625 414520 345646
rect 414478 247616 414534 247625
rect 414478 247551 414534 247560
rect 414584 235414 414612 345918
rect 414572 235408 414624 235414
rect 414572 235350 414624 235356
rect 414676 147286 414704 457234
rect 414756 457156 414808 457162
rect 414756 457098 414808 457104
rect 414768 149666 414796 457098
rect 414848 457020 414900 457026
rect 414848 456962 414900 456968
rect 414756 149660 414808 149666
rect 414756 149602 414808 149608
rect 414860 149530 414888 456962
rect 414940 455864 414992 455870
rect 414940 455806 414992 455812
rect 414848 149524 414900 149530
rect 414848 149466 414900 149472
rect 414952 149161 414980 455806
rect 415032 454980 415084 454986
rect 415032 454922 415084 454928
rect 415044 149598 415072 454922
rect 415214 451616 415270 451625
rect 415214 451551 415270 451560
rect 415122 449984 415178 449993
rect 415122 449919 415178 449928
rect 415032 149592 415084 149598
rect 415032 149534 415084 149540
rect 414938 149152 414994 149161
rect 414938 149087 414994 149096
rect 415136 147422 415164 449919
rect 415228 158166 415256 451551
rect 415320 249014 415348 458458
rect 415858 452024 415914 452033
rect 415858 451959 415914 451968
rect 415872 346361 415900 451959
rect 415858 346352 415914 346361
rect 415858 346287 415914 346296
rect 415860 345908 415912 345914
rect 415860 345850 415912 345856
rect 415872 340202 415900 345850
rect 415952 345840 416004 345846
rect 415952 345782 416004 345788
rect 415964 345574 415992 345782
rect 415952 345568 416004 345574
rect 415952 345510 416004 345516
rect 415860 340196 415912 340202
rect 415860 340138 415912 340144
rect 415308 249008 415360 249014
rect 415308 248950 415360 248956
rect 415860 237448 415912 237454
rect 415860 237390 415912 237396
rect 415676 234796 415728 234802
rect 415676 234738 415728 234744
rect 415216 158160 415268 158166
rect 415216 158102 415268 158108
rect 415124 147416 415176 147422
rect 415124 147358 415176 147364
rect 414664 147280 414716 147286
rect 414664 147222 414716 147228
rect 415688 146130 415716 234738
rect 415768 234728 415820 234734
rect 415768 234670 415820 234676
rect 415780 146266 415808 234670
rect 415872 149734 415900 237390
rect 415964 235346 415992 345510
rect 415952 235340 416004 235346
rect 415952 235282 416004 235288
rect 415860 149728 415912 149734
rect 415860 149670 415912 149676
rect 415768 146260 415820 146266
rect 415768 146202 415820 146208
rect 415676 146124 415728 146130
rect 415676 146066 415728 146072
rect 416056 48278 416084 462334
rect 416136 457632 416188 457638
rect 416136 457574 416188 457580
rect 416148 49230 416176 457574
rect 416320 456272 416372 456278
rect 416320 456214 416372 456220
rect 416228 455456 416280 455462
rect 416228 455398 416280 455404
rect 416136 49224 416188 49230
rect 416136 49166 416188 49172
rect 416044 48272 416096 48278
rect 416044 48214 416096 48220
rect 416240 47297 416268 455398
rect 416332 347410 416360 456214
rect 417516 453620 417568 453626
rect 417516 453562 417568 453568
rect 416964 452736 417016 452742
rect 416964 452678 417016 452684
rect 416594 451888 416650 451897
rect 416594 451823 416650 451832
rect 416410 451752 416466 451761
rect 416410 451687 416466 451696
rect 416320 347404 416372 347410
rect 416320 347346 416372 347352
rect 416320 345636 416372 345642
rect 416320 345578 416372 345584
rect 416332 235550 416360 345578
rect 416320 235544 416372 235550
rect 416320 235486 416372 235492
rect 416332 234666 416360 235486
rect 416320 234660 416372 234666
rect 416320 234602 416372 234608
rect 416320 146260 416372 146266
rect 416320 146202 416372 146208
rect 416226 47288 416282 47297
rect 416226 47223 416282 47232
rect 416332 45558 416360 146202
rect 416424 47161 416452 451687
rect 416504 451512 416556 451518
rect 416504 451454 416556 451460
rect 416516 346934 416544 451454
rect 416504 346928 416556 346934
rect 416504 346870 416556 346876
rect 416504 340196 416556 340202
rect 416504 340138 416556 340144
rect 416516 235686 416544 340138
rect 416504 235680 416556 235686
rect 416504 235622 416556 235628
rect 416516 234802 416544 235622
rect 416504 234796 416556 234802
rect 416504 234738 416556 234744
rect 416504 234660 416556 234666
rect 416504 234602 416556 234608
rect 416516 145926 416544 234602
rect 416504 145920 416556 145926
rect 416504 145862 416556 145868
rect 416410 47152 416466 47161
rect 416410 47087 416466 47096
rect 416320 45552 416372 45558
rect 416320 45494 416372 45500
rect 416516 45286 416544 145862
rect 416608 49026 416636 451823
rect 416688 449676 416740 449682
rect 416688 449618 416740 449624
rect 416700 349246 416728 449618
rect 416780 382968 416832 382974
rect 416780 382910 416832 382916
rect 416792 382809 416820 382910
rect 416778 382800 416834 382809
rect 416778 382735 416834 382744
rect 416872 381540 416924 381546
rect 416872 381482 416924 381488
rect 416884 381041 416912 381482
rect 416870 381032 416926 381041
rect 416870 380967 416926 380976
rect 416780 380180 416832 380186
rect 416780 380122 416832 380128
rect 416792 379953 416820 380122
rect 416778 379944 416834 379953
rect 416778 379879 416834 379888
rect 416780 378820 416832 378826
rect 416780 378762 416832 378768
rect 416792 378185 416820 378762
rect 416778 378176 416834 378185
rect 416778 378111 416834 378120
rect 416976 358057 417004 452678
rect 417424 451444 417476 451450
rect 417424 451386 417476 451392
rect 417330 386880 417386 386889
rect 417330 386815 417386 386824
rect 417238 386336 417294 386345
rect 417238 386271 417294 386280
rect 417252 385937 417280 386271
rect 417238 385928 417294 385937
rect 417238 385863 417294 385872
rect 417146 358320 417202 358329
rect 417146 358255 417202 358264
rect 416962 358048 417018 358057
rect 416962 357983 417018 357992
rect 416688 349240 416740 349246
rect 416688 349182 416740 349188
rect 416688 345840 416740 345846
rect 416688 345782 416740 345788
rect 416700 345506 416728 345782
rect 416688 345500 416740 345506
rect 416688 345442 416740 345448
rect 416700 235754 416728 345442
rect 417054 285696 417110 285705
rect 417054 285631 417110 285640
rect 416870 281072 416926 281081
rect 416870 281007 416926 281016
rect 416688 235748 416740 235754
rect 416688 235690 416740 235696
rect 416700 234734 416728 235690
rect 416688 234728 416740 234734
rect 416688 234670 416740 234676
rect 416884 182073 416912 281007
rect 417068 186017 417096 285631
rect 417160 258126 417188 358255
rect 417252 285977 417280 385863
rect 417344 286929 417372 386815
rect 417436 347750 417464 451386
rect 417528 383654 417556 453562
rect 417700 452872 417752 452878
rect 417700 452814 417752 452820
rect 417608 452804 417660 452810
rect 417608 452746 417660 452752
rect 417620 386345 417648 452746
rect 417712 386889 417740 452814
rect 417698 386880 417754 386889
rect 417698 386815 417754 386824
rect 417606 386336 417662 386345
rect 417606 386271 417662 386280
rect 417882 383752 417938 383761
rect 417882 383687 417938 383696
rect 417896 383654 417924 383687
rect 417528 383626 417924 383654
rect 417514 382800 417570 382809
rect 417514 382735 417570 382744
rect 417424 347744 417476 347750
rect 417424 347686 417476 347692
rect 417528 287054 417556 382735
rect 417790 381032 417846 381041
rect 417790 380967 417846 380976
rect 417698 379944 417754 379953
rect 417698 379879 417754 379888
rect 417606 378176 417662 378185
rect 417606 378111 417662 378120
rect 417436 287026 417556 287054
rect 417330 286920 417386 286929
rect 417330 286855 417386 286864
rect 417238 285968 417294 285977
rect 417238 285903 417294 285912
rect 417252 285705 417280 285903
rect 417238 285696 417294 285705
rect 417238 285631 417294 285640
rect 417238 283792 417294 283801
rect 417238 283727 417294 283736
rect 417148 258120 417200 258126
rect 417148 258062 417200 258068
rect 417148 235340 417200 235346
rect 417148 235282 417200 235288
rect 417054 186008 417110 186017
rect 417054 185943 417110 185952
rect 416870 182064 416926 182073
rect 416870 181999 416926 182008
rect 416688 146124 416740 146130
rect 416688 146066 416740 146072
rect 416596 49020 416648 49026
rect 416596 48962 416648 48968
rect 416700 45490 416728 146066
rect 417068 85921 417096 185943
rect 417160 146266 417188 235282
rect 417252 183841 417280 283727
rect 417344 186969 417372 286855
rect 417436 282849 417464 287026
rect 417422 282840 417478 282849
rect 417422 282775 417478 282784
rect 417330 186960 417386 186969
rect 417330 186895 417386 186904
rect 417238 183832 417294 183841
rect 417238 183767 417294 183776
rect 417436 182889 417464 282775
rect 417620 278769 417648 378111
rect 417712 279993 417740 379879
rect 417804 281081 417832 380967
rect 417896 283801 417924 383626
rect 418080 358329 418108 508263
rect 418816 500274 418844 700266
rect 462332 587178 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 479524 700324 479576 700330
rect 479524 700266 479576 700272
rect 462320 587172 462372 587178
rect 462320 587114 462372 587120
rect 479536 585818 479564 700266
rect 479524 585812 479576 585818
rect 479524 585754 479576 585760
rect 494072 584458 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 542372 588606 542400 702406
rect 559668 699718 559696 703520
rect 558184 699712 558236 699718
rect 558184 699654 558236 699660
rect 559656 699712 559708 699718
rect 559656 699654 559708 699660
rect 542360 588600 542412 588606
rect 542360 588542 542412 588548
rect 551008 585200 551060 585206
rect 551006 585168 551008 585177
rect 557540 585200 557592 585206
rect 551060 585168 551062 585177
rect 557540 585142 557592 585148
rect 551006 585103 551062 585112
rect 494060 584452 494112 584458
rect 494060 584394 494112 584400
rect 418804 500268 418856 500274
rect 418804 500210 418856 500216
rect 557552 498234 557580 585142
rect 551928 498228 551980 498234
rect 551928 498170 551980 498176
rect 557540 498228 557592 498234
rect 557540 498170 557592 498176
rect 441618 498128 441674 498137
rect 441618 498063 441674 498072
rect 444378 498128 444434 498137
rect 444378 498063 444434 498072
rect 448518 498128 448574 498137
rect 448518 498063 448574 498072
rect 451278 498128 451334 498137
rect 451278 498063 451334 498072
rect 454682 498128 454738 498137
rect 454682 498063 454738 498072
rect 473358 498128 473414 498137
rect 480350 498128 480406 498137
rect 473358 498063 473414 498072
rect 476764 498092 476816 498098
rect 436190 497312 436246 497321
rect 436190 497247 436246 497256
rect 436098 497176 436154 497185
rect 436204 497146 436232 497247
rect 436098 497111 436154 497120
rect 436192 497140 436244 497146
rect 436112 497078 436140 497111
rect 436192 497082 436244 497088
rect 436100 497072 436152 497078
rect 436100 497014 436152 497020
rect 437478 496904 437534 496913
rect 437478 496839 437534 496848
rect 438858 496904 438914 496913
rect 438858 496839 438914 496848
rect 440238 496904 440294 496913
rect 440238 496839 440294 496848
rect 437492 494766 437520 496839
rect 437480 494760 437532 494766
rect 437480 494702 437532 494708
rect 438872 483682 438900 496839
rect 438860 483676 438912 483682
rect 438860 483618 438912 483624
rect 418896 459808 418948 459814
rect 418896 459750 418948 459756
rect 418804 458312 418856 458318
rect 418804 458254 418856 458260
rect 418066 358320 418122 358329
rect 418066 358255 418122 358264
rect 418160 349920 418212 349926
rect 418160 349862 418212 349868
rect 418172 349654 418200 349862
rect 418160 349648 418212 349654
rect 418160 349590 418212 349596
rect 418068 349036 418120 349042
rect 418068 348978 418120 348984
rect 418080 347818 418108 348978
rect 418712 348696 418764 348702
rect 418712 348638 418764 348644
rect 418724 347954 418752 348638
rect 418712 347948 418764 347954
rect 418712 347890 418764 347896
rect 418068 347812 418120 347818
rect 418068 347754 418120 347760
rect 417976 347744 418028 347750
rect 417976 347686 418028 347692
rect 417988 347070 418016 347686
rect 417976 347064 418028 347070
rect 417976 347006 418028 347012
rect 417882 283792 417938 283801
rect 417882 283727 417938 283736
rect 417790 281072 417846 281081
rect 417790 281007 417846 281016
rect 417698 279984 417754 279993
rect 417698 279919 417754 279928
rect 417606 278760 417662 278769
rect 417606 278695 417662 278704
rect 417712 258074 417740 279919
rect 417884 259412 417936 259418
rect 417884 259354 417936 259360
rect 417896 258097 417924 259354
rect 417528 258046 417740 258074
rect 417882 258088 417938 258097
rect 417422 182880 417478 182889
rect 417422 182815 417478 182824
rect 417238 182064 417294 182073
rect 417238 181999 417294 182008
rect 417252 181121 417280 181999
rect 417238 181112 417294 181121
rect 417238 181047 417294 181056
rect 417148 146260 417200 146266
rect 417148 146202 417200 146208
rect 417054 85912 417110 85921
rect 417054 85847 417110 85856
rect 417252 81025 417280 181047
rect 417332 134428 417384 134434
rect 417332 134370 417384 134376
rect 417238 81016 417294 81025
rect 417238 80951 417294 80960
rect 416780 59356 416832 59362
rect 416780 59298 416832 59304
rect 416792 58041 416820 59298
rect 416778 58032 416834 58041
rect 416778 57967 416834 57976
rect 417344 48006 417372 134370
rect 417436 82929 417464 182815
rect 417528 180033 417556 258046
rect 417882 258023 417938 258032
rect 417700 253224 417752 253230
rect 417700 253166 417752 253172
rect 417712 235958 417740 253166
rect 417790 247616 417846 247625
rect 417790 247551 417846 247560
rect 417700 235952 417752 235958
rect 417700 235894 417752 235900
rect 417514 180024 417570 180033
rect 417514 179959 417570 179968
rect 417528 179489 417556 179959
rect 417514 179480 417570 179489
rect 417514 179415 417570 179424
rect 417712 161474 417740 235894
rect 417620 161446 417740 161474
rect 417620 158409 417648 161446
rect 417606 158400 417662 158409
rect 417606 158335 417662 158344
rect 417422 82920 417478 82929
rect 417422 82855 417478 82864
rect 417620 58313 417648 158335
rect 417700 158160 417752 158166
rect 417698 158128 417700 158137
rect 417752 158128 417754 158137
rect 417698 158063 417754 158072
rect 417700 149728 417752 149734
rect 417700 149670 417752 149676
rect 417606 58304 417662 58313
rect 417606 58239 417662 58248
rect 417712 49910 417740 149670
rect 417804 146985 417832 247551
rect 417988 235278 418016 347006
rect 418080 235890 418108 347754
rect 418618 346352 418674 346361
rect 418618 346287 418674 346296
rect 418632 345681 418660 346287
rect 418618 345672 418674 345681
rect 418618 345607 418674 345616
rect 418632 342990 418660 345607
rect 418620 342984 418672 342990
rect 418620 342926 418672 342932
rect 418618 258360 418674 258369
rect 418618 258295 418674 258304
rect 418632 258126 418660 258295
rect 418620 258120 418672 258126
rect 418620 258062 418672 258068
rect 418632 253230 418660 258062
rect 418620 253224 418672 253230
rect 418620 253166 418672 253172
rect 418342 249520 418398 249529
rect 418342 249455 418398 249464
rect 418068 235884 418120 235890
rect 418068 235826 418120 235832
rect 417976 235272 418028 235278
rect 417976 235214 418028 235220
rect 417882 186960 417938 186969
rect 417882 186895 417938 186904
rect 417790 146976 417846 146985
rect 417790 146911 417846 146920
rect 417792 146260 417844 146266
rect 417792 146202 417844 146208
rect 417804 145858 417832 146202
rect 417792 145852 417844 145858
rect 417792 145794 417844 145800
rect 417700 49904 417752 49910
rect 417700 49846 417752 49852
rect 417332 48000 417384 48006
rect 417332 47942 417384 47948
rect 417804 46442 417832 145794
rect 417896 86873 417924 186895
rect 417974 183832 418030 183841
rect 417974 183767 418030 183776
rect 417882 86864 417938 86873
rect 417882 86799 417938 86808
rect 417988 83745 418016 183767
rect 418080 147121 418108 235826
rect 418356 147354 418384 249455
rect 418724 248414 418752 347890
rect 418816 248878 418844 458254
rect 418908 348514 418936 459750
rect 440252 457502 440280 496839
rect 441632 486470 441660 498063
rect 442998 497040 443054 497049
rect 442998 496975 443054 496984
rect 441620 486464 441672 486470
rect 441620 486406 441672 486412
rect 443012 461650 443040 496975
rect 443090 496904 443146 496913
rect 443090 496839 443146 496848
rect 443104 487830 443132 496839
rect 443092 487824 443144 487830
rect 443092 487766 443144 487772
rect 443000 461644 443052 461650
rect 443000 461586 443052 461592
rect 444392 458862 444420 498063
rect 447138 497040 447194 497049
rect 447138 496975 447194 496984
rect 445758 496904 445814 496913
rect 445758 496839 445814 496848
rect 445772 464370 445800 496839
rect 445760 464364 445812 464370
rect 445760 464306 445812 464312
rect 447152 463010 447180 496975
rect 447230 496904 447286 496913
rect 447230 496839 447286 496848
rect 447244 468586 447272 496839
rect 448532 496194 448560 498063
rect 449990 497040 450046 497049
rect 449990 496975 450046 496984
rect 449898 496904 449954 496913
rect 449898 496839 449954 496848
rect 448520 496188 448572 496194
rect 448520 496130 448572 496136
rect 449912 469946 449940 496839
rect 450004 472666 450032 496975
rect 449992 472660 450044 472666
rect 449992 472602 450044 472608
rect 449900 469940 449952 469946
rect 449900 469882 449952 469888
rect 447232 468580 447284 468586
rect 447232 468522 447284 468528
rect 447140 463004 447192 463010
rect 447140 462946 447192 462952
rect 451292 460290 451320 498063
rect 452658 497584 452714 497593
rect 452658 497519 452714 497528
rect 452672 497214 452700 497519
rect 452660 497208 452712 497214
rect 452660 497150 452712 497156
rect 451370 496904 451426 496913
rect 451370 496839 451426 496848
rect 452750 496904 452806 496913
rect 452750 496839 452806 496848
rect 454038 496904 454094 496913
rect 454038 496839 454094 496848
rect 451384 471306 451412 496839
rect 452764 474094 452792 496839
rect 454052 493338 454080 496839
rect 454040 493332 454092 493338
rect 454040 493274 454092 493280
rect 454696 475386 454724 498063
rect 455418 497176 455474 497185
rect 455418 497111 455474 497120
rect 455432 496126 455460 497111
rect 473372 497078 473400 498063
rect 480350 498063 480352 498072
rect 476764 498034 476816 498040
rect 480404 498063 480406 498072
rect 480352 498034 480404 498040
rect 457444 497072 457496 497078
rect 456890 497040 456946 497049
rect 473360 497072 473412 497078
rect 457444 497014 457496 497020
rect 458270 497040 458326 497049
rect 456890 496975 456946 496984
rect 456798 496904 456854 496913
rect 456798 496839 456854 496848
rect 455420 496120 455472 496126
rect 455420 496062 455472 496068
rect 456812 489258 456840 496839
rect 456904 490618 456932 496975
rect 456892 490612 456944 490618
rect 456892 490554 456944 490560
rect 456800 489252 456852 489258
rect 456800 489194 456852 489200
rect 454684 475380 454736 475386
rect 454684 475322 454736 475328
rect 452752 474088 452804 474094
rect 452752 474030 452804 474036
rect 451372 471300 451424 471306
rect 451372 471242 451424 471248
rect 457456 468518 457484 497014
rect 458270 496975 458326 496984
rect 459558 497040 459614 497049
rect 470782 497040 470838 497049
rect 459558 496975 459560 496984
rect 458178 496904 458234 496913
rect 458178 496839 458234 496848
rect 458192 476814 458220 496839
rect 458284 491978 458312 496975
rect 459612 496975 459614 496984
rect 464344 497004 464396 497010
rect 459560 496946 459612 496952
rect 473360 497014 473412 497020
rect 476118 497040 476174 497049
rect 470782 496975 470838 496984
rect 476118 496975 476120 496984
rect 464344 496946 464396 496952
rect 460938 496904 460994 496913
rect 460938 496839 460994 496848
rect 462318 496904 462374 496913
rect 462318 496839 462374 496848
rect 458272 491972 458324 491978
rect 458272 491914 458324 491920
rect 460952 479602 460980 496839
rect 460940 479596 460992 479602
rect 460940 479538 460992 479544
rect 462332 478174 462360 496839
rect 462320 478168 462372 478174
rect 462320 478110 462372 478116
rect 458180 476808 458232 476814
rect 458180 476750 458232 476756
rect 464356 469878 464384 496946
rect 470796 496942 470824 496975
rect 476172 496975 476174 496984
rect 476120 496946 476172 496952
rect 470784 496936 470836 496942
rect 465078 496904 465134 496913
rect 465078 496839 465134 496848
rect 467838 496904 467894 496913
rect 470784 496878 470836 496884
rect 475384 496936 475436 496942
rect 475384 496878 475436 496884
rect 467838 496839 467894 496848
rect 472624 496868 472676 496874
rect 465092 481030 465120 496839
rect 467852 482322 467880 496839
rect 472624 496810 472676 496816
rect 467840 482316 467892 482322
rect 467840 482258 467892 482264
rect 465080 481024 465132 481030
rect 465080 480966 465132 480972
rect 464344 469872 464396 469878
rect 464344 469814 464396 469820
rect 457444 468512 457496 468518
rect 457444 468454 457496 468460
rect 472636 465798 472664 496810
rect 475396 467158 475424 496878
rect 475384 467152 475436 467158
rect 475384 467094 475436 467100
rect 472624 465792 472676 465798
rect 472624 465734 472676 465740
rect 451280 460284 451332 460290
rect 451280 460226 451332 460232
rect 476776 460222 476804 498034
rect 485778 497992 485834 498001
rect 485778 497927 485834 497936
rect 485792 497282 485820 497927
rect 485780 497276 485832 497282
rect 485780 497218 485832 497224
rect 483018 497176 483074 497185
rect 483018 497111 483074 497120
rect 483032 496942 483060 497111
rect 483020 496936 483072 496942
rect 477498 496904 477554 496913
rect 483020 496878 483072 496884
rect 477498 496839 477500 496848
rect 477552 496839 477554 496848
rect 477500 496810 477552 496816
rect 476764 460216 476816 460222
rect 476764 460158 476816 460164
rect 493416 459604 493468 459610
rect 493416 459546 493468 459552
rect 444380 458856 444432 458862
rect 444380 458798 444432 458804
rect 493428 458182 493456 459546
rect 493416 458176 493468 458182
rect 493416 458118 493468 458124
rect 440240 457496 440292 457502
rect 440240 457438 440292 457444
rect 419264 457224 419316 457230
rect 419264 457166 419316 457172
rect 418988 454504 419040 454510
rect 418988 454446 419040 454452
rect 419000 348770 419028 454446
rect 419080 451308 419132 451314
rect 419080 451250 419132 451256
rect 418988 348764 419040 348770
rect 418988 348706 419040 348712
rect 419092 348702 419120 451250
rect 419080 348696 419132 348702
rect 419080 348638 419132 348644
rect 418908 348486 419120 348514
rect 418896 347404 418948 347410
rect 418896 347346 418948 347352
rect 418908 346458 418936 347346
rect 419092 347206 419120 348486
rect 419276 347274 419304 457166
rect 419356 456204 419408 456210
rect 419356 456146 419408 456152
rect 419368 347410 419396 456146
rect 419630 452704 419686 452713
rect 419630 452639 419686 452648
rect 419448 349648 419500 349654
rect 419448 349590 419500 349596
rect 419356 347404 419408 347410
rect 419356 347346 419408 347352
rect 419172 347268 419224 347274
rect 419172 347210 419224 347216
rect 419264 347268 419316 347274
rect 419264 347210 419316 347216
rect 419080 347200 419132 347206
rect 419080 347142 419132 347148
rect 418896 346452 418948 346458
rect 418896 346394 418948 346400
rect 418908 345014 418936 346394
rect 418908 344986 419028 345014
rect 418896 342984 418948 342990
rect 418896 342926 418948 342932
rect 418804 248872 418856 248878
rect 418804 248814 418856 248820
rect 418540 248386 418752 248414
rect 418540 247722 418568 248386
rect 418528 247716 418580 247722
rect 418528 247658 418580 247664
rect 418436 234660 418488 234666
rect 418436 234602 418488 234608
rect 418344 147348 418396 147354
rect 418344 147290 418396 147296
rect 418066 147112 418122 147121
rect 418066 147047 418122 147056
rect 418448 147014 418476 234602
rect 418436 147008 418488 147014
rect 418436 146950 418488 146956
rect 418540 135250 418568 247658
rect 418620 243568 418672 243574
rect 418620 243510 418672 243516
rect 418632 235521 418660 243510
rect 418908 238754 418936 342926
rect 419000 243574 419028 344986
rect 418988 243568 419040 243574
rect 418988 243510 419040 243516
rect 418908 238726 419028 238754
rect 419000 235929 419028 238726
rect 418986 235920 419042 235929
rect 418986 235855 419042 235864
rect 418618 235512 418674 235521
rect 419092 235482 419120 347142
rect 419184 346594 419212 347210
rect 419172 346588 419224 346594
rect 419172 346530 419224 346536
rect 419184 235657 419212 346530
rect 419170 235648 419226 235657
rect 419170 235583 419226 235592
rect 418618 235447 418674 235456
rect 419080 235476 419132 235482
rect 418632 146878 418660 235447
rect 419080 235418 419132 235424
rect 418988 235408 419040 235414
rect 418988 235350 419040 235356
rect 418712 235136 418764 235142
rect 418712 235078 418764 235084
rect 418724 147218 418752 235078
rect 418896 235068 418948 235074
rect 418896 235010 418948 235016
rect 418712 147212 418764 147218
rect 418712 147154 418764 147160
rect 418710 147112 418766 147121
rect 418710 147047 418766 147056
rect 418620 146872 418672 146878
rect 418620 146814 418672 146820
rect 418528 135244 418580 135250
rect 418528 135186 418580 135192
rect 418540 134434 418568 135186
rect 418528 134428 418580 134434
rect 418528 134370 418580 134376
rect 417974 83736 418030 83745
rect 417974 83671 418030 83680
rect 418724 49978 418752 147047
rect 418802 146976 418858 146985
rect 418802 146911 418858 146920
rect 418712 49972 418764 49978
rect 418712 49914 418764 49920
rect 418816 48822 418844 146911
rect 418908 146810 418936 235010
rect 418896 146804 418948 146810
rect 418896 146746 418948 146752
rect 418804 48816 418856 48822
rect 418804 48758 418856 48764
rect 418908 47598 418936 146746
rect 419000 145790 419028 235350
rect 419092 234666 419120 235418
rect 419080 234660 419132 234666
rect 419080 234602 419132 234608
rect 419184 171134 419212 235583
rect 419276 235074 419304 347210
rect 419368 235142 419396 347346
rect 419460 235618 419488 349590
rect 419540 349104 419592 349110
rect 419540 349046 419592 349052
rect 419552 347886 419580 349046
rect 419540 347880 419592 347886
rect 419538 347848 419540 347857
rect 419592 347848 419594 347857
rect 419538 347783 419594 347792
rect 419644 347313 419672 452639
rect 419998 449848 420054 449857
rect 419998 449783 420054 449792
rect 420012 348838 420040 449783
rect 551940 435402 551968 498170
rect 558196 465730 558224 699654
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 558918 578640 558974 578649
rect 558918 578575 558974 578584
rect 558276 510672 558328 510678
rect 558276 510614 558328 510620
rect 558288 498846 558316 510614
rect 558276 498840 558328 498846
rect 558276 498782 558328 498788
rect 558184 465724 558236 465730
rect 558184 465666 558236 465672
rect 558276 461168 558328 461174
rect 558276 461110 558328 461116
rect 558182 456240 558238 456249
rect 558182 456175 558238 456184
rect 551928 435396 551980 435402
rect 551928 435338 551980 435344
rect 557540 435396 557592 435402
rect 557540 435338 557592 435344
rect 557552 433537 557580 435338
rect 557538 433528 557594 433537
rect 557538 433463 557594 433472
rect 478510 349888 478566 349897
rect 478510 349823 478566 349832
rect 483478 349888 483534 349897
rect 483478 349823 483534 349832
rect 485962 349888 486018 349897
rect 485962 349823 486018 349832
rect 492586 349888 492642 349897
rect 492586 349823 492588 349832
rect 452566 349752 452622 349761
rect 452566 349687 452622 349696
rect 452580 349654 452608 349687
rect 452568 349648 452620 349654
rect 452568 349590 452620 349596
rect 420000 348832 420052 348838
rect 420000 348774 420052 348780
rect 436098 347712 436154 347721
rect 436098 347647 436154 347656
rect 437018 347712 437074 347721
rect 437018 347647 437074 347656
rect 438030 347712 438086 347721
rect 438030 347647 438086 347656
rect 439594 347712 439650 347721
rect 439594 347647 439650 347656
rect 440514 347712 440570 347721
rect 440514 347647 440570 347656
rect 441618 347712 441674 347721
rect 441618 347647 441674 347656
rect 443090 347712 443146 347721
rect 443090 347647 443146 347656
rect 444194 347712 444250 347721
rect 444194 347647 444250 347656
rect 445298 347712 445354 347721
rect 445298 347647 445354 347656
rect 446402 347712 446458 347721
rect 446402 347647 446458 347656
rect 447138 347712 447194 347721
rect 447138 347647 447194 347656
rect 448242 347712 448298 347721
rect 448242 347647 448298 347656
rect 448518 347712 448574 347721
rect 448518 347647 448574 347656
rect 449898 347712 449954 347721
rect 449898 347647 449954 347656
rect 450634 347712 450690 347721
rect 450634 347647 450690 347656
rect 451370 347712 451426 347721
rect 451370 347647 451426 347656
rect 419724 347336 419776 347342
rect 419630 347304 419686 347313
rect 419724 347278 419776 347284
rect 419630 347239 419686 347248
rect 419632 347132 419684 347138
rect 419632 347074 419684 347080
rect 419644 346866 419672 347074
rect 419632 346860 419684 346866
rect 419632 346802 419684 346808
rect 419644 238746 419672 346802
rect 419736 346526 419764 347278
rect 436112 347274 436140 347647
rect 437032 347410 437060 347647
rect 437020 347404 437072 347410
rect 437020 347346 437072 347352
rect 436744 347336 436796 347342
rect 436744 347278 436796 347284
rect 436100 347268 436152 347274
rect 436100 347210 436152 347216
rect 419816 347132 419868 347138
rect 419816 347074 419868 347080
rect 419828 346934 419856 347074
rect 419816 346928 419868 346934
rect 419814 346896 419816 346905
rect 419868 346896 419870 346905
rect 419814 346831 419870 346840
rect 419724 346520 419776 346526
rect 419724 346462 419776 346468
rect 419736 248414 419764 346462
rect 420000 346112 420052 346118
rect 420000 346054 420052 346060
rect 419908 345772 419960 345778
rect 419908 345714 419960 345720
rect 419736 248386 419856 248414
rect 419632 238740 419684 238746
rect 419632 238682 419684 238688
rect 419644 237454 419672 238682
rect 419828 238678 419856 248386
rect 419816 238672 419868 238678
rect 419816 238614 419868 238620
rect 419632 237448 419684 237454
rect 419632 237390 419684 237396
rect 419448 235612 419500 235618
rect 419448 235554 419500 235560
rect 419356 235136 419408 235142
rect 419356 235078 419408 235084
rect 419264 235068 419316 235074
rect 419264 235010 419316 235016
rect 419184 171106 419396 171134
rect 419080 147212 419132 147218
rect 419080 147154 419132 147160
rect 418988 145784 419040 145790
rect 418988 145726 419040 145732
rect 418896 47592 418948 47598
rect 418896 47534 418948 47540
rect 419000 46510 419028 145726
rect 419092 47530 419120 147154
rect 419368 147150 419396 171106
rect 419356 147144 419408 147150
rect 419356 147086 419408 147092
rect 419264 147008 419316 147014
rect 419264 146950 419316 146956
rect 419172 146872 419224 146878
rect 419172 146814 419224 146820
rect 419184 47666 419212 146814
rect 419276 47870 419304 146950
rect 419264 47864 419316 47870
rect 419264 47806 419316 47812
rect 419368 47734 419396 147086
rect 419460 146130 419488 235554
rect 419540 235272 419592 235278
rect 419540 235214 419592 235220
rect 419448 146124 419500 146130
rect 419448 146066 419500 146072
rect 419356 47728 419408 47734
rect 419356 47670 419408 47676
rect 419172 47660 419224 47666
rect 419172 47602 419224 47608
rect 419080 47524 419132 47530
rect 419080 47466 419132 47472
rect 418988 46504 419040 46510
rect 418988 46446 419040 46452
rect 417792 46436 417844 46442
rect 417792 46378 417844 46384
rect 416688 45484 416740 45490
rect 416688 45426 416740 45432
rect 419460 45422 419488 146066
rect 419552 145994 419580 235214
rect 419724 235204 419776 235210
rect 419724 235146 419776 235152
rect 419736 151814 419764 235146
rect 419644 151786 419764 151814
rect 419644 147082 419672 151786
rect 419632 147076 419684 147082
rect 419632 147018 419684 147024
rect 419540 145988 419592 145994
rect 419540 145930 419592 145936
rect 419644 47802 419672 147018
rect 419724 146940 419776 146946
rect 419724 146882 419776 146888
rect 419736 47938 419764 146882
rect 419828 146198 419856 238614
rect 419920 235822 419948 345714
rect 420012 345506 420040 346054
rect 436756 345506 436784 347278
rect 438044 346458 438072 347647
rect 439608 346594 439636 347647
rect 440528 347138 440556 347647
rect 440516 347132 440568 347138
rect 440516 347074 440568 347080
rect 439596 346588 439648 346594
rect 439596 346530 439648 346536
rect 441632 346458 441660 347647
rect 443104 347342 443132 347647
rect 443092 347336 443144 347342
rect 443092 347278 443144 347284
rect 444208 347138 444236 347647
rect 444196 347132 444248 347138
rect 444196 347074 444248 347080
rect 445312 346594 445340 347647
rect 446416 346662 446444 347647
rect 447152 346730 447180 347647
rect 448256 347478 448284 347647
rect 448244 347472 448296 347478
rect 448244 347414 448296 347420
rect 448532 346798 448560 347647
rect 448520 346792 448572 346798
rect 448520 346734 448572 346740
rect 447140 346724 447192 346730
rect 447140 346666 447192 346672
rect 446404 346656 446456 346662
rect 446404 346598 446456 346604
rect 445300 346588 445352 346594
rect 445300 346530 445352 346536
rect 438032 346452 438084 346458
rect 438032 346394 438084 346400
rect 438860 346452 438912 346458
rect 438860 346394 438912 346400
rect 441620 346452 441672 346458
rect 441620 346394 441672 346400
rect 438872 345681 438900 346394
rect 438858 345672 438914 345681
rect 438858 345607 438914 345616
rect 445312 345574 445340 346530
rect 446416 345982 446444 346598
rect 446404 345976 446456 345982
rect 446404 345918 446456 345924
rect 447152 345642 447180 346666
rect 448532 345914 448560 346734
rect 449912 346458 449940 347647
rect 450648 347546 450676 347647
rect 450636 347540 450688 347546
rect 450636 347482 450688 347488
rect 451384 347070 451412 347647
rect 452580 347546 452608 349590
rect 478524 349586 478552 349823
rect 478512 349580 478564 349586
rect 478512 349522 478564 349528
rect 483492 349518 483520 349823
rect 483480 349512 483532 349518
rect 483480 349454 483532 349460
rect 485976 349450 486004 349823
rect 492640 349823 492642 349832
rect 492588 349794 492640 349800
rect 488262 349752 488318 349761
rect 488262 349687 488318 349696
rect 491022 349752 491078 349761
rect 491022 349687 491078 349696
rect 508502 349752 508558 349761
rect 508502 349687 508558 349696
rect 520922 349752 520978 349761
rect 520922 349687 520978 349696
rect 485964 349444 486016 349450
rect 485964 349386 486016 349392
rect 488276 349382 488304 349687
rect 488264 349376 488316 349382
rect 488264 349318 488316 349324
rect 491036 349314 491064 349687
rect 505926 349616 505982 349625
rect 505926 349551 505982 349560
rect 491024 349308 491076 349314
rect 491024 349250 491076 349256
rect 498474 349072 498530 349081
rect 498474 349007 498530 349016
rect 500958 349072 501014 349081
rect 500958 349007 501014 349016
rect 503442 349072 503498 349081
rect 503442 349007 503498 349016
rect 498488 348634 498516 349007
rect 500972 348838 501000 349007
rect 500960 348832 501012 348838
rect 500960 348774 501012 348780
rect 498476 348628 498528 348634
rect 498476 348570 498528 348576
rect 503456 348498 503484 349007
rect 505940 348770 505968 349551
rect 508516 349178 508544 349687
rect 515862 349616 515918 349625
rect 515862 349551 515918 349560
rect 508504 349172 508556 349178
rect 508504 349114 508556 349120
rect 510986 349072 511042 349081
rect 510986 349007 511042 349016
rect 505928 348764 505980 348770
rect 505928 348706 505980 348712
rect 503444 348492 503496 348498
rect 503444 348434 503496 348440
rect 511000 348430 511028 349007
rect 515876 348702 515904 349551
rect 520936 349246 520964 349687
rect 520924 349240 520976 349246
rect 520924 349182 520976 349188
rect 523314 349072 523370 349081
rect 523314 349007 523370 349016
rect 515864 348696 515916 348702
rect 515864 348638 515916 348644
rect 523328 348566 523356 349007
rect 523316 348560 523368 348566
rect 523316 348502 523368 348508
rect 510988 348424 511040 348430
rect 510988 348366 511040 348372
rect 455788 347948 455840 347954
rect 455788 347890 455840 347896
rect 455800 347721 455828 347890
rect 458180 347880 458232 347886
rect 458180 347822 458232 347828
rect 456984 347812 457036 347818
rect 456984 347754 457036 347760
rect 456996 347721 457024 347754
rect 458192 347750 458220 347822
rect 462228 347812 462280 347818
rect 462228 347754 462280 347760
rect 458180 347744 458232 347750
rect 453026 347712 453082 347721
rect 453026 347647 453082 347656
rect 453578 347712 453634 347721
rect 453578 347647 453634 347656
rect 455234 347712 455290 347721
rect 455234 347647 455290 347656
rect 455786 347712 455842 347721
rect 455786 347647 455842 347656
rect 456154 347712 456210 347721
rect 456154 347647 456210 347656
rect 456982 347712 457038 347721
rect 456982 347647 457038 347656
rect 458086 347712 458142 347721
rect 459468 347744 459520 347750
rect 458180 347686 458232 347692
rect 458362 347712 458418 347721
rect 458086 347647 458142 347656
rect 458362 347647 458364 347656
rect 452568 347540 452620 347546
rect 452568 347482 452620 347488
rect 452568 347268 452620 347274
rect 452568 347210 452620 347216
rect 452580 347070 452608 347210
rect 453040 347070 453068 347647
rect 453592 347614 453620 347647
rect 453580 347608 453632 347614
rect 453580 347550 453632 347556
rect 451372 347064 451424 347070
rect 451372 347006 451424 347012
rect 452568 347064 452620 347070
rect 452568 347006 452620 347012
rect 453028 347064 453080 347070
rect 453028 347006 453080 347012
rect 453040 346526 453068 347006
rect 455248 346526 455276 347647
rect 455800 347614 455828 347647
rect 455788 347608 455840 347614
rect 455788 347550 455840 347556
rect 456168 347002 456196 347647
rect 458100 347206 458128 347647
rect 458416 347647 458418 347656
rect 459466 347712 459468 347721
rect 459520 347712 459522 347721
rect 459466 347647 459522 347656
rect 460938 347712 460994 347721
rect 460938 347647 460994 347656
rect 461490 347712 461546 347721
rect 462240 347682 462268 347754
rect 478052 347744 478104 347750
rect 462778 347712 462834 347721
rect 461490 347647 461546 347656
rect 462228 347676 462280 347682
rect 458364 347618 458416 347624
rect 456800 347200 456852 347206
rect 456800 347142 456852 347148
rect 458088 347200 458140 347206
rect 458088 347142 458140 347148
rect 456156 346996 456208 347002
rect 456156 346938 456208 346944
rect 456812 346866 456840 347142
rect 460570 347032 460626 347041
rect 460570 346967 460626 346976
rect 456800 346860 456852 346866
rect 456800 346802 456852 346808
rect 453028 346520 453080 346526
rect 453028 346462 453080 346468
rect 455236 346520 455288 346526
rect 455236 346462 455288 346468
rect 449900 346452 449952 346458
rect 449900 346394 449952 346400
rect 448520 345908 448572 345914
rect 448520 345850 448572 345856
rect 449912 345846 449940 346394
rect 449900 345840 449952 345846
rect 449900 345782 449952 345788
rect 455248 345778 455276 346462
rect 460584 346118 460612 346967
rect 459560 346112 459612 346118
rect 459560 346054 459612 346060
rect 460572 346112 460624 346118
rect 460572 346054 460624 346060
rect 455236 345772 455288 345778
rect 455236 345714 455288 345720
rect 459572 345710 459600 346054
rect 460952 346050 460980 347647
rect 461504 347342 461532 347647
rect 462778 347647 462834 347656
rect 463514 347712 463570 347721
rect 463514 347647 463570 347656
rect 463882 347712 463938 347721
rect 463882 347647 463938 347656
rect 465170 347712 465226 347721
rect 465170 347647 465226 347656
rect 465722 347712 465778 347721
rect 465722 347647 465778 347656
rect 467378 347712 467434 347721
rect 467378 347647 467434 347656
rect 468666 347712 468722 347721
rect 468666 347647 468722 347656
rect 469770 347712 469826 347721
rect 469770 347647 469826 347656
rect 471242 347712 471298 347721
rect 471242 347647 471298 347656
rect 472070 347712 472126 347721
rect 472070 347647 472126 347656
rect 473358 347712 473414 347721
rect 473358 347647 473414 347656
rect 474370 347712 474426 347721
rect 474370 347647 474426 347656
rect 475658 347712 475714 347721
rect 475658 347647 475660 347656
rect 462228 347618 462280 347624
rect 461492 347336 461544 347342
rect 461492 347278 461544 347284
rect 462792 347138 462820 347647
rect 462780 347132 462832 347138
rect 462780 347074 462832 347080
rect 460940 346044 460992 346050
rect 460940 345986 460992 345992
rect 459560 345704 459612 345710
rect 459560 345646 459612 345652
rect 447140 345636 447192 345642
rect 447140 345578 447192 345584
rect 445300 345568 445352 345574
rect 445300 345510 445352 345516
rect 420000 345500 420052 345506
rect 420000 345442 420052 345448
rect 436744 345500 436796 345506
rect 436744 345442 436796 345448
rect 419908 235816 419960 235822
rect 419908 235758 419960 235764
rect 419920 146946 419948 235758
rect 420012 235210 420040 345442
rect 463528 345370 463556 347647
rect 463896 346594 463924 347647
rect 465184 346662 465212 347647
rect 465262 347032 465318 347041
rect 465262 346967 465318 346976
rect 465172 346656 465224 346662
rect 465172 346598 465224 346604
rect 463884 346588 463936 346594
rect 463884 346530 463936 346536
rect 465276 346186 465304 346967
rect 465736 346730 465764 347647
rect 467392 346798 467420 347647
rect 467930 347576 467986 347585
rect 467930 347511 467986 347520
rect 467380 346792 467432 346798
rect 467380 346734 467432 346740
rect 465724 346724 465776 346730
rect 465724 346666 465776 346672
rect 465264 346180 465316 346186
rect 465264 346122 465316 346128
rect 463516 345364 463568 345370
rect 463516 345306 463568 345312
rect 467944 345030 467972 347511
rect 468680 346458 468708 347647
rect 469784 347274 469812 347647
rect 471256 347546 471284 347647
rect 471244 347540 471296 347546
rect 471244 347482 471296 347488
rect 469772 347268 469824 347274
rect 469772 347210 469824 347216
rect 472084 347070 472112 347647
rect 472072 347064 472124 347070
rect 472072 347006 472124 347012
rect 473372 346526 473400 347647
rect 474384 347614 474412 347647
rect 475712 347647 475714 347656
rect 476946 347712 477002 347721
rect 478050 347712 478052 347721
rect 478104 347712 478106 347721
rect 476946 347647 477002 347656
rect 477408 347676 477460 347682
rect 475660 347618 475712 347624
rect 474372 347608 474424 347614
rect 474372 347550 474424 347556
rect 476960 347206 476988 347647
rect 478050 347647 478106 347656
rect 479154 347712 479210 347721
rect 479154 347647 479156 347656
rect 477408 347618 477460 347624
rect 479208 347647 479210 347656
rect 513378 347712 513434 347721
rect 513378 347647 513434 347656
rect 518346 347712 518402 347721
rect 518346 347647 518402 347656
rect 525890 347712 525946 347721
rect 525890 347647 525946 347656
rect 479156 347618 479208 347624
rect 476948 347200 477000 347206
rect 476948 347142 477000 347148
rect 473360 346520 473412 346526
rect 473360 346462 473412 346468
rect 468668 346452 468720 346458
rect 468668 346394 468720 346400
rect 477420 346118 477448 347618
rect 513392 346254 513420 347647
rect 518360 346322 518388 347647
rect 525904 346390 525932 347647
rect 525892 346384 525944 346390
rect 525892 346326 525944 346332
rect 518348 346316 518400 346322
rect 518348 346258 518400 346264
rect 513380 346248 513432 346254
rect 513380 346190 513432 346196
rect 477408 346112 477460 346118
rect 477408 346054 477460 346060
rect 467932 345024 467984 345030
rect 467932 344966 467984 344972
rect 557552 335510 557580 433463
rect 558196 353258 558224 456175
rect 558288 431934 558316 461110
rect 558276 431928 558328 431934
rect 558276 431870 558328 431876
rect 558932 429729 558960 578575
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 562324 563100 562376 563106
rect 562324 563042 562376 563048
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 562336 489190 562364 563042
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 563704 536852 563756 536858
rect 563704 536794 563756 536800
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 562324 489184 562376 489190
rect 562324 489126 562376 489132
rect 563716 474026 563744 536794
rect 580170 524512 580226 524521
rect 565084 524476 565136 524482
rect 580170 524447 580172 524456
rect 565084 524418 565136 524424
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 565096 479534 565124 524418
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580276 480962 580304 577623
rect 580264 480956 580316 480962
rect 580264 480898 580316 480904
rect 565084 479528 565136 479534
rect 565084 479470 565136 479476
rect 563704 474020 563756 474026
rect 563704 473962 563756 473968
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 577688 466880 577740 466886
rect 577688 466822 577740 466828
rect 577504 466540 577556 466546
rect 577504 466482 577556 466488
rect 559564 461236 559616 461242
rect 559564 461178 559616 461184
rect 558918 429720 558974 429729
rect 558918 429655 558974 429664
rect 558184 353252 558236 353258
rect 558184 353194 558236 353200
rect 551008 335504 551060 335510
rect 551006 335472 551008 335481
rect 557540 335504 557592 335510
rect 551060 335472 551062 335481
rect 557540 335446 557592 335452
rect 551006 335407 551062 335416
rect 485962 249792 486018 249801
rect 485962 249727 485964 249736
rect 486016 249727 486018 249736
rect 488262 249792 488318 249801
rect 488262 249727 488318 249736
rect 491022 249792 491078 249801
rect 491022 249727 491078 249736
rect 495898 249792 495954 249801
rect 495898 249727 495954 249736
rect 498474 249792 498530 249801
rect 498474 249727 498530 249736
rect 500958 249792 501014 249801
rect 500958 249727 501014 249736
rect 503534 249792 503590 249801
rect 503534 249727 503590 249736
rect 485964 249698 486016 249704
rect 488276 249694 488304 249727
rect 488264 249688 488316 249694
rect 470966 249656 471022 249665
rect 470966 249591 471022 249600
rect 483478 249656 483534 249665
rect 488264 249630 488316 249636
rect 491036 249626 491064 249727
rect 483478 249591 483534 249600
rect 491024 249620 491076 249626
rect 470980 248946 471008 249591
rect 473634 249384 473690 249393
rect 473634 249319 473690 249328
rect 470968 248940 471020 248946
rect 470968 248882 471020 248888
rect 473648 248878 473676 249319
rect 483492 249014 483520 249591
rect 491024 249562 491076 249568
rect 495912 249558 495940 249727
rect 495900 249552 495952 249558
rect 495900 249494 495952 249500
rect 498488 249490 498516 249727
rect 498476 249484 498528 249490
rect 498476 249426 498528 249432
rect 500972 249422 501000 249727
rect 500960 249416 501012 249422
rect 500960 249358 501012 249364
rect 503548 249354 503576 249727
rect 505926 249656 505982 249665
rect 505926 249591 505982 249600
rect 508502 249656 508558 249665
rect 508502 249591 508558 249600
rect 515862 249656 515918 249665
rect 515862 249591 515918 249600
rect 520922 249656 520978 249665
rect 520922 249591 520978 249600
rect 503536 249348 503588 249354
rect 503536 249290 503588 249296
rect 505940 249286 505968 249591
rect 505928 249280 505980 249286
rect 505928 249222 505980 249228
rect 508516 249218 508544 249591
rect 508504 249212 508556 249218
rect 508504 249154 508556 249160
rect 515876 249150 515904 249591
rect 515864 249144 515916 249150
rect 515864 249086 515916 249092
rect 520936 249082 520964 249591
rect 520924 249076 520976 249082
rect 520924 249018 520976 249024
rect 483480 249008 483532 249014
rect 483480 248950 483532 248956
rect 473636 248872 473688 248878
rect 473636 248814 473688 248820
rect 455420 248328 455472 248334
rect 443182 248296 443238 248305
rect 443182 248231 443238 248240
rect 447138 248296 447194 248305
rect 447138 248231 447194 248240
rect 449806 248296 449862 248305
rect 450174 248296 450230 248305
rect 449862 248254 449940 248282
rect 449806 248231 449862 248240
rect 443196 247994 443224 248231
rect 447152 248130 447180 248231
rect 447140 248124 447192 248130
rect 447140 248066 447192 248072
rect 444472 248056 444524 248062
rect 444472 247998 444524 248004
rect 443184 247988 443236 247994
rect 443184 247930 443236 247936
rect 444196 247988 444248 247994
rect 444196 247930 444248 247936
rect 436098 247344 436154 247353
rect 436098 247279 436154 247288
rect 420000 235204 420052 235210
rect 420000 235146 420052 235152
rect 436112 235142 436140 247279
rect 436190 247072 436246 247081
rect 436190 247007 436246 247016
rect 437478 247072 437534 247081
rect 437478 247007 437534 247016
rect 438858 247072 438914 247081
rect 438858 247007 438914 247016
rect 440238 247072 440294 247081
rect 440238 247007 440294 247016
rect 441618 247072 441674 247081
rect 441618 247007 441674 247016
rect 436100 235136 436152 235142
rect 436100 235078 436152 235084
rect 436204 235074 436232 247007
rect 437492 235521 437520 247007
rect 438872 235657 438900 247007
rect 440252 235793 440280 247007
rect 441632 235929 441660 247007
rect 444208 246922 444236 247930
rect 444286 247072 444342 247081
rect 444484 247058 444512 247998
rect 447140 247920 447192 247926
rect 447140 247862 447192 247868
rect 445760 247376 445812 247382
rect 445760 247318 445812 247324
rect 444342 247030 444512 247058
rect 444286 247007 444342 247016
rect 444208 246894 444420 246922
rect 441618 235920 441674 235929
rect 441618 235855 441674 235864
rect 440238 235784 440294 235793
rect 440238 235719 440294 235728
rect 438858 235648 438914 235657
rect 438858 235583 438914 235592
rect 437478 235512 437534 235521
rect 437478 235447 437534 235456
rect 444392 235210 444420 246894
rect 444484 235482 444512 247030
rect 445666 247072 445722 247081
rect 445772 247058 445800 247318
rect 445722 247030 445800 247058
rect 445666 247007 445722 247016
rect 444472 235476 444524 235482
rect 444472 235418 444524 235424
rect 445772 235346 445800 247030
rect 447046 247072 447102 247081
rect 447152 247058 447180 247862
rect 449912 247654 449940 248254
rect 450174 248231 450230 248240
rect 450358 248296 450414 248305
rect 450358 248231 450414 248240
rect 451370 248296 451426 248305
rect 451370 248231 451426 248240
rect 452658 248296 452714 248305
rect 452658 248231 452660 248240
rect 450188 248130 450216 248231
rect 450372 248198 450400 248231
rect 450360 248192 450412 248198
rect 450360 248134 450412 248140
rect 450176 248124 450228 248130
rect 450176 248066 450228 248072
rect 451280 248124 451332 248130
rect 451280 248066 451332 248072
rect 449900 247648 449952 247654
rect 449900 247590 449952 247596
rect 448520 247580 448572 247586
rect 448520 247522 448572 247528
rect 447102 247030 447180 247058
rect 447046 247007 447102 247016
rect 447152 235414 447180 247030
rect 448426 247072 448482 247081
rect 448532 247058 448560 247522
rect 448482 247030 448560 247058
rect 448426 247007 448482 247016
rect 448532 235550 448560 247030
rect 449912 235686 449940 247590
rect 451292 235754 451320 248066
rect 451384 247858 451412 248231
rect 452712 248231 452714 248240
rect 455418 248296 455420 248305
rect 455472 248296 455474 248305
rect 455418 248231 455474 248240
rect 462318 248296 462374 248305
rect 462318 248231 462374 248240
rect 467838 248296 467894 248305
rect 467838 248231 467894 248240
rect 452660 248202 452712 248208
rect 462332 248062 462360 248231
rect 467852 248130 467880 248231
rect 467840 248124 467892 248130
rect 467840 248066 467892 248072
rect 462320 248056 462372 248062
rect 460938 248024 460994 248033
rect 460938 247959 460994 247968
rect 461122 248024 461178 248033
rect 462320 247998 462372 248004
rect 465078 248024 465134 248033
rect 461122 247959 461124 247968
rect 460952 247874 460980 247959
rect 461176 247959 461178 247968
rect 465078 247959 465134 247968
rect 461124 247930 461176 247936
rect 465092 247926 465120 247959
rect 465080 247920 465132 247926
rect 461122 247888 461178 247897
rect 451372 247852 451424 247858
rect 451372 247794 451424 247800
rect 452476 247852 452528 247858
rect 460952 247846 461122 247874
rect 461122 247823 461178 247832
rect 463698 247888 463754 247897
rect 465080 247862 465132 247868
rect 469218 247888 469274 247897
rect 463698 247823 463754 247832
rect 469218 247823 469220 247832
rect 452476 247794 452528 247800
rect 452488 246922 452516 247794
rect 455880 247784 455932 247790
rect 455880 247726 455932 247732
rect 455892 247625 455920 247726
rect 462228 247716 462280 247722
rect 462228 247658 462280 247664
rect 462240 247625 462268 247658
rect 455878 247616 455934 247625
rect 455878 247551 455934 247560
rect 462226 247616 462282 247625
rect 462226 247551 462282 247560
rect 452752 247512 452804 247518
rect 452752 247454 452804 247460
rect 457994 247480 458050 247489
rect 452566 247072 452622 247081
rect 452764 247058 452792 247454
rect 457994 247415 458050 247424
rect 458272 247444 458324 247450
rect 455420 247240 455472 247246
rect 455420 247182 455472 247188
rect 454040 247172 454092 247178
rect 454040 247114 454092 247120
rect 452622 247030 452792 247058
rect 452566 247007 452622 247016
rect 452488 246894 452700 246922
rect 451280 235748 451332 235754
rect 451280 235690 451332 235696
rect 449900 235680 449952 235686
rect 449900 235622 449952 235628
rect 448520 235544 448572 235550
rect 448520 235486 448572 235492
rect 447140 235408 447192 235414
rect 447140 235350 447192 235356
rect 445760 235340 445812 235346
rect 445760 235282 445812 235288
rect 452672 235278 452700 246894
rect 452764 235618 452792 247030
rect 453946 247072 454002 247081
rect 454052 247058 454080 247114
rect 454002 247030 454080 247058
rect 453946 247007 454002 247016
rect 454052 238678 454080 247030
rect 455326 247072 455382 247081
rect 455432 247058 455460 247182
rect 455382 247030 455460 247058
rect 455326 247007 455382 247016
rect 454040 238672 454092 238678
rect 454040 238614 454092 238620
rect 455432 235822 455460 247030
rect 458008 246922 458036 247415
rect 458272 247386 458324 247392
rect 458086 247072 458142 247081
rect 458284 247058 458312 247386
rect 463712 247382 463740 247823
rect 469272 247823 469274 247832
rect 473358 247888 473414 247897
rect 473358 247823 473414 247832
rect 469220 247794 469272 247800
rect 473372 247790 473400 247823
rect 473360 247784 473412 247790
rect 466458 247752 466514 247761
rect 473360 247726 473412 247732
rect 478878 247752 478934 247761
rect 466458 247687 466514 247696
rect 478878 247687 478880 247696
rect 466472 247654 466500 247687
rect 478932 247687 478934 247696
rect 478880 247658 478932 247664
rect 466460 247648 466512 247654
rect 465078 247616 465134 247625
rect 466460 247590 466512 247596
rect 470782 247616 470838 247625
rect 465078 247551 465080 247560
rect 465132 247551 465134 247560
rect 470782 247551 470838 247560
rect 465080 247522 465132 247528
rect 470796 247518 470824 247551
rect 470784 247512 470836 247518
rect 470784 247454 470836 247460
rect 476118 247480 476174 247489
rect 476118 247415 476120 247424
rect 476172 247415 476174 247424
rect 476120 247386 476172 247392
rect 463700 247376 463752 247382
rect 459466 247344 459522 247353
rect 459522 247314 459600 247330
rect 463700 247318 463752 247324
rect 471978 247344 472034 247353
rect 459522 247308 459612 247314
rect 459522 247302 459560 247308
rect 459466 247279 459522 247288
rect 471978 247279 472034 247288
rect 473358 247344 473414 247353
rect 473358 247279 473414 247288
rect 477498 247344 477554 247353
rect 477498 247279 477500 247288
rect 459560 247250 459612 247256
rect 458142 247030 458312 247058
rect 458086 247007 458142 247016
rect 458008 246894 458220 246922
rect 458192 235890 458220 246894
rect 458284 238746 458312 247030
rect 458272 238740 458324 238746
rect 458272 238682 458324 238688
rect 459572 238649 459600 247250
rect 471992 247178 472020 247279
rect 473372 247246 473400 247279
rect 477552 247279 477554 247288
rect 477500 247250 477552 247256
rect 473360 247240 473412 247246
rect 473360 247182 473412 247188
rect 471980 247172 472032 247178
rect 471980 247114 472032 247120
rect 480534 247072 480590 247081
rect 480534 247007 480590 247016
rect 492678 247072 492734 247081
rect 492678 247007 492734 247016
rect 510618 247072 510674 247081
rect 510618 247007 510674 247016
rect 513378 247072 513434 247081
rect 513378 247007 513434 247016
rect 523038 247072 523094 247081
rect 523038 247007 523094 247016
rect 525798 247072 525854 247081
rect 525798 247007 525800 247016
rect 480548 245478 480576 247007
rect 492692 245546 492720 247007
rect 510632 246906 510660 247007
rect 513392 246974 513420 247007
rect 513380 246968 513432 246974
rect 513380 246910 513432 246916
rect 510620 246900 510672 246906
rect 510620 246842 510672 246848
rect 523052 245614 523080 247007
rect 525852 247007 525854 247016
rect 525800 246978 525852 246984
rect 523040 245608 523092 245614
rect 523040 245550 523092 245556
rect 492680 245540 492732 245546
rect 492680 245482 492732 245488
rect 480536 245472 480588 245478
rect 480536 245414 480588 245420
rect 459558 238640 459614 238649
rect 459558 238575 459614 238584
rect 550824 235952 550876 235958
rect 550824 235894 550876 235900
rect 557448 235952 557500 235958
rect 557552 235906 557580 335446
rect 558932 329225 558960 429655
rect 559576 419490 559604 461178
rect 563704 461100 563756 461106
rect 563704 461042 563756 461048
rect 559564 419484 559616 419490
rect 559564 419426 559616 419432
rect 558918 329216 558974 329225
rect 558918 329151 558974 329160
rect 558184 246424 558236 246430
rect 558184 246366 558236 246372
rect 557632 240780 557684 240786
rect 557632 240722 557684 240728
rect 557500 235900 557580 235906
rect 557448 235894 557580 235900
rect 458180 235884 458232 235890
rect 458180 235826 458232 235832
rect 455420 235816 455472 235822
rect 455420 235758 455472 235764
rect 452752 235612 452804 235618
rect 452752 235554 452804 235560
rect 452660 235272 452712 235278
rect 452660 235214 452712 235220
rect 444380 235204 444432 235210
rect 444380 235146 444432 235152
rect 550836 235113 550864 235894
rect 557460 235878 557580 235894
rect 550822 235104 550878 235113
rect 436192 235068 436244 235074
rect 550822 235039 550878 235048
rect 436192 235010 436244 235016
rect 557552 234598 557580 235878
rect 556804 234592 556856 234598
rect 556804 234534 556856 234540
rect 557540 234592 557592 234598
rect 557540 234534 557592 234540
rect 458086 149832 458142 149841
rect 458086 149767 458142 149776
rect 478510 149832 478566 149841
rect 478510 149767 478566 149776
rect 480902 149832 480958 149841
rect 480902 149767 480958 149776
rect 483478 149832 483534 149841
rect 483478 149767 483534 149776
rect 485962 149832 486018 149841
rect 485962 149767 486018 149776
rect 458100 149734 458128 149767
rect 458088 149728 458140 149734
rect 440054 149696 440110 149705
rect 458088 149670 458140 149676
rect 440054 149631 440110 149640
rect 438214 149560 438270 149569
rect 438214 149495 438270 149504
rect 436098 147656 436154 147665
rect 436098 147591 436154 147600
rect 437018 147656 437074 147665
rect 437018 147591 437074 147600
rect 437938 147656 437994 147665
rect 437938 147591 437994 147600
rect 419908 146940 419960 146946
rect 419908 146882 419960 146888
rect 430578 146840 430634 146849
rect 436112 146810 436140 147591
rect 437032 147218 437060 147591
rect 437020 147212 437072 147218
rect 437020 147154 437072 147160
rect 437952 146878 437980 147591
rect 437940 146872 437992 146878
rect 437940 146814 437992 146820
rect 430578 146775 430634 146784
rect 436100 146804 436152 146810
rect 430592 146742 430620 146775
rect 436100 146746 436152 146752
rect 438228 146742 438256 149495
rect 439594 147656 439650 147665
rect 439594 147591 439650 147600
rect 439608 147150 439636 147591
rect 440068 147257 440096 149631
rect 456798 149560 456854 149569
rect 456798 149495 456854 149504
rect 443090 147656 443146 147665
rect 443090 147591 443146 147600
rect 444194 147656 444250 147665
rect 444194 147591 444250 147600
rect 445298 147656 445354 147665
rect 445298 147591 445354 147600
rect 446402 147656 446458 147665
rect 446402 147591 446458 147600
rect 447138 147656 447194 147665
rect 447138 147591 447194 147600
rect 448242 147656 448298 147665
rect 448242 147591 448298 147600
rect 448518 147656 448574 147665
rect 448518 147591 448574 147600
rect 449898 147656 449954 147665
rect 449898 147591 449954 147600
rect 450634 147656 450690 147665
rect 450634 147591 450690 147600
rect 451278 147656 451334 147665
rect 451278 147591 451334 147600
rect 452566 147656 452622 147665
rect 452566 147591 452622 147600
rect 453394 147656 453450 147665
rect 453394 147591 453450 147600
rect 453578 147656 453634 147665
rect 453578 147591 453634 147600
rect 454590 147656 454646 147665
rect 454590 147591 454646 147600
rect 455970 147656 456026 147665
rect 455970 147591 456026 147600
rect 440240 147280 440292 147286
rect 440054 147248 440110 147257
rect 440054 147183 440110 147192
rect 440238 147248 440240 147257
rect 440292 147248 440294 147257
rect 440238 147183 440294 147192
rect 439596 147144 439648 147150
rect 439596 147086 439648 147092
rect 443104 147082 443132 147591
rect 443092 147076 443144 147082
rect 443092 147018 443144 147024
rect 444208 147014 444236 147591
rect 444196 147008 444248 147014
rect 444196 146950 444248 146956
rect 445312 146878 445340 147591
rect 445300 146872 445352 146878
rect 445300 146814 445352 146820
rect 430580 146736 430632 146742
rect 430580 146678 430632 146684
rect 438216 146736 438268 146742
rect 438216 146678 438268 146684
rect 419816 146192 419868 146198
rect 419816 146134 419868 146140
rect 419724 47932 419776 47938
rect 419724 47874 419776 47880
rect 419632 47796 419684 47802
rect 419632 47738 419684 47744
rect 419828 46578 419856 146134
rect 420000 145988 420052 145994
rect 420000 145930 420052 145936
rect 419816 46572 419868 46578
rect 419816 46514 419868 46520
rect 419448 45416 419500 45422
rect 419448 45358 419500 45364
rect 420012 45354 420040 145930
rect 445312 145858 445340 146814
rect 446416 146470 446444 147591
rect 447152 146810 447180 147591
rect 448256 147422 448284 147591
rect 448244 147416 448296 147422
rect 448244 147358 448296 147364
rect 447140 146804 447192 146810
rect 447140 146746 447192 146752
rect 446404 146464 446456 146470
rect 446404 146406 446456 146412
rect 445300 145852 445352 145858
rect 445300 145794 445352 145800
rect 446416 145790 446444 146406
rect 447152 145926 447180 146746
rect 448532 146742 448560 147591
rect 448520 146736 448572 146742
rect 448520 146678 448572 146684
rect 448532 146062 448560 146678
rect 449912 146674 449940 147591
rect 450648 147354 450676 147591
rect 450636 147348 450688 147354
rect 450636 147290 450688 147296
rect 449900 146668 449952 146674
rect 449900 146610 449952 146616
rect 449912 146266 449940 146610
rect 449900 146260 449952 146266
rect 449900 146202 449952 146208
rect 448520 146056 448572 146062
rect 448520 145998 448572 146004
rect 451292 145994 451320 147591
rect 452476 146600 452528 146606
rect 452476 146542 452528 146548
rect 452488 145994 452516 146542
rect 452580 146538 452608 147591
rect 452568 146532 452620 146538
rect 452568 146474 452620 146480
rect 452580 146130 452608 146474
rect 453408 146198 453436 147591
rect 453592 147490 453620 147591
rect 453580 147484 453632 147490
rect 453580 147426 453632 147432
rect 454604 146946 454632 147591
rect 455984 147558 456012 147591
rect 455972 147552 456024 147558
rect 455972 147494 456024 147500
rect 454592 146940 454644 146946
rect 454592 146882 454644 146888
rect 456812 146334 456840 149495
rect 458100 147558 458128 149670
rect 478524 149666 478552 149767
rect 478512 149660 478564 149666
rect 478512 149602 478564 149608
rect 480916 149598 480944 149767
rect 480904 149592 480956 149598
rect 463514 149560 463570 149569
rect 463514 149495 463570 149504
rect 465998 149560 466054 149569
rect 465998 149495 466054 149504
rect 468298 149560 468354 149569
rect 468298 149495 468354 149504
rect 470966 149560 471022 149569
rect 480904 149534 480956 149540
rect 483492 149530 483520 149767
rect 470966 149495 471022 149504
rect 483480 149524 483532 149530
rect 459466 148744 459522 148753
rect 459466 148679 459522 148688
rect 459480 148345 459508 148679
rect 459466 148336 459522 148345
rect 459466 148271 459522 148280
rect 458362 147656 458418 147665
rect 459480 147626 459508 148271
rect 463528 148238 463556 149495
rect 466012 148306 466040 149495
rect 468312 149054 468340 149495
rect 468300 149048 468352 149054
rect 468300 148990 468352 148996
rect 470980 148986 471008 149495
rect 483480 149466 483532 149472
rect 485976 149462 486004 149767
rect 488262 149696 488318 149705
rect 488262 149631 488318 149640
rect 491022 149696 491078 149705
rect 491022 149631 491078 149640
rect 495898 149696 495954 149705
rect 495898 149631 495954 149640
rect 503534 149696 503590 149705
rect 503534 149631 503590 149640
rect 485964 149456 486016 149462
rect 485964 149398 486016 149404
rect 488276 149394 488304 149631
rect 488264 149388 488316 149394
rect 488264 149330 488316 149336
rect 491036 149326 491064 149631
rect 491024 149320 491076 149326
rect 491024 149262 491076 149268
rect 495912 149258 495940 149631
rect 495900 149252 495952 149258
rect 495900 149194 495952 149200
rect 503548 149190 503576 149631
rect 505926 149560 505982 149569
rect 505926 149495 505982 149504
rect 508502 149560 508558 149569
rect 508502 149495 508558 149504
rect 510986 149560 511042 149569
rect 510986 149495 511042 149504
rect 515862 149560 515918 149569
rect 515862 149495 515918 149504
rect 518438 149560 518494 149569
rect 518438 149495 518494 149504
rect 503536 149184 503588 149190
rect 503536 149126 503588 149132
rect 470968 148980 471020 148986
rect 470968 148922 471020 148928
rect 505940 148918 505968 149495
rect 505928 148912 505980 148918
rect 505928 148854 505980 148860
rect 508516 148850 508544 149495
rect 508504 148844 508556 148850
rect 508504 148786 508556 148792
rect 511000 148782 511028 149495
rect 513378 149016 513434 149025
rect 513378 148951 513434 148960
rect 510988 148776 511040 148782
rect 510988 148718 511040 148724
rect 513392 148714 513420 148951
rect 513380 148708 513432 148714
rect 513380 148650 513432 148656
rect 515876 148646 515904 149495
rect 518452 149122 518480 149495
rect 518440 149116 518492 149122
rect 518440 149058 518492 149064
rect 520922 149016 520978 149025
rect 520922 148951 520978 148960
rect 523314 149016 523370 149025
rect 523314 148951 523370 148960
rect 525890 149016 525946 149025
rect 525890 148951 525946 148960
rect 515864 148640 515916 148646
rect 515864 148582 515916 148588
rect 520936 148578 520964 148951
rect 520924 148572 520976 148578
rect 520924 148514 520976 148520
rect 523328 148510 523356 148951
rect 523316 148504 523368 148510
rect 523316 148446 523368 148452
rect 525904 148442 525932 148951
rect 525892 148436 525944 148442
rect 525892 148378 525944 148384
rect 531044 148368 531096 148374
rect 531044 148310 531096 148316
rect 466000 148300 466052 148306
rect 466000 148242 466052 148248
rect 463516 148232 463568 148238
rect 463516 148174 463568 148180
rect 461674 147656 461730 147665
rect 458362 147591 458364 147600
rect 458416 147591 458418 147600
rect 459468 147620 459520 147626
rect 458364 147562 458416 147568
rect 461674 147591 461730 147600
rect 462778 147656 462834 147665
rect 462778 147591 462834 147600
rect 463882 147656 463938 147665
rect 463882 147591 463938 147600
rect 465170 147656 465226 147665
rect 465170 147591 465226 147600
rect 466274 147656 466330 147665
rect 466274 147591 466330 147600
rect 467562 147656 467618 147665
rect 467562 147591 467618 147600
rect 468666 147656 468722 147665
rect 468666 147591 468722 147600
rect 469770 147656 469826 147665
rect 469770 147591 469826 147600
rect 471058 147656 471114 147665
rect 471058 147591 471114 147600
rect 472162 147656 472218 147665
rect 472162 147591 472218 147600
rect 473358 147656 473414 147665
rect 473358 147591 473414 147600
rect 474094 147656 474150 147665
rect 474094 147591 474150 147600
rect 476946 147656 477002 147665
rect 476946 147591 477002 147600
rect 478050 147656 478106 147665
rect 478050 147591 478052 147600
rect 459468 147562 459520 147568
rect 458088 147552 458140 147558
rect 458088 147494 458140 147500
rect 461688 147082 461716 147591
rect 461676 147076 461728 147082
rect 461676 147018 461728 147024
rect 462792 147014 462820 147591
rect 462780 147008 462832 147014
rect 462780 146950 462832 146956
rect 463896 146878 463924 147591
rect 463884 146872 463936 146878
rect 463884 146814 463936 146820
rect 465184 146470 465212 147591
rect 466288 146810 466316 147591
rect 466276 146804 466328 146810
rect 466276 146746 466328 146752
rect 467576 146742 467604 147591
rect 467564 146736 467616 146742
rect 467564 146678 467616 146684
rect 468680 146674 468708 147591
rect 468668 146668 468720 146674
rect 468668 146610 468720 146616
rect 469784 146606 469812 147591
rect 469772 146600 469824 146606
rect 469772 146542 469824 146548
rect 471072 146538 471100 147591
rect 471060 146532 471112 146538
rect 471060 146474 471112 146480
rect 465172 146464 465224 146470
rect 465172 146406 465224 146412
rect 472176 146402 472204 147591
rect 473372 146946 473400 147591
rect 473360 146940 473412 146946
rect 473360 146882 473412 146888
rect 472164 146396 472216 146402
rect 472164 146338 472216 146344
rect 474108 146334 474136 147591
rect 476960 147558 476988 147591
rect 478104 147591 478106 147600
rect 478052 147562 478104 147568
rect 476948 147552 477000 147558
rect 476948 147494 477000 147500
rect 456800 146328 456852 146334
rect 456800 146270 456852 146276
rect 474096 146328 474148 146334
rect 474096 146270 474148 146276
rect 453396 146192 453448 146198
rect 453396 146134 453448 146140
rect 452568 146124 452620 146130
rect 452568 146066 452620 146072
rect 451280 145988 451332 145994
rect 451280 145930 451332 145936
rect 452476 145988 452528 145994
rect 452476 145930 452528 145936
rect 447140 145920 447192 145926
rect 447140 145862 447192 145868
rect 446404 145784 446456 145790
rect 446404 145726 446456 145732
rect 456812 135250 456840 146270
rect 531056 144906 531084 148310
rect 531044 144900 531096 144906
rect 531044 144842 531096 144848
rect 536840 144900 536892 144906
rect 536840 144842 536892 144848
rect 536852 138718 536880 144842
rect 536840 138712 536892 138718
rect 536840 138654 536892 138660
rect 556816 136610 556844 234534
rect 557644 229265 557672 240722
rect 557630 229256 557686 229265
rect 557630 229191 557686 229200
rect 556896 138712 556948 138718
rect 556896 138654 556948 138660
rect 551928 136604 551980 136610
rect 551928 136546 551980 136552
rect 556804 136604 556856 136610
rect 556804 136546 556856 136552
rect 551940 136513 551968 136546
rect 551926 136504 551982 136513
rect 551926 136439 551982 136448
rect 456800 135244 456852 135250
rect 456800 135186 456852 135192
rect 556908 110430 556936 138654
rect 556896 110424 556948 110430
rect 556896 110366 556948 110372
rect 456984 49972 457036 49978
rect 456984 49914 457036 49920
rect 456996 49881 457024 49914
rect 458088 49904 458140 49910
rect 456982 49872 457038 49881
rect 456982 49807 457038 49816
rect 458086 49872 458088 49881
rect 458140 49872 458142 49881
rect 458086 49807 458142 49816
rect 478510 49872 478566 49881
rect 478510 49807 478512 49816
rect 436098 48240 436154 48249
rect 436098 48175 436154 48184
rect 437018 48240 437074 48249
rect 437018 48175 437074 48184
rect 438122 48240 438178 48249
rect 438122 48175 438178 48184
rect 439594 48240 439650 48249
rect 439594 48175 439650 48184
rect 443090 48240 443146 48249
rect 443090 48175 443146 48184
rect 444286 48240 444342 48249
rect 444286 48175 444342 48184
rect 448242 48240 448298 48249
rect 448242 48175 448244 48184
rect 436112 47598 436140 48175
rect 436100 47592 436152 47598
rect 436100 47534 436152 47540
rect 437032 47530 437060 48175
rect 438136 47666 438164 48175
rect 439608 47734 439636 48175
rect 443104 47734 443132 48175
rect 444300 47870 444328 48175
rect 448296 48175 448298 48184
rect 450634 48240 450690 48249
rect 450634 48175 450690 48184
rect 453578 48240 453634 48249
rect 453578 48175 453634 48184
rect 454590 48240 454646 48249
rect 454590 48175 454646 48184
rect 455878 48240 455934 48249
rect 455878 48175 455934 48184
rect 448244 48146 448296 48152
rect 445298 48104 445354 48113
rect 445298 48039 445354 48048
rect 446402 48104 446458 48113
rect 446402 48039 446458 48048
rect 449530 48104 449586 48113
rect 450648 48074 450676 48175
rect 453592 48142 453620 48175
rect 453580 48136 453632 48142
rect 452290 48104 452346 48113
rect 449530 48039 449586 48048
rect 450636 48068 450688 48074
rect 444288 47864 444340 47870
rect 444288 47806 444340 47812
rect 439596 47728 439648 47734
rect 439596 47670 439648 47676
rect 443092 47728 443144 47734
rect 443092 47670 443144 47676
rect 444300 47666 444328 47806
rect 438124 47660 438176 47666
rect 438124 47602 438176 47608
rect 444288 47660 444340 47666
rect 444288 47602 444340 47608
rect 437020 47524 437072 47530
rect 437020 47466 437072 47472
rect 445312 47122 445340 48039
rect 445300 47116 445352 47122
rect 445300 47058 445352 47064
rect 445312 46442 445340 47058
rect 446416 47054 446444 48039
rect 447506 47560 447562 47569
rect 447506 47495 447562 47504
rect 447520 47258 447548 47495
rect 449544 47394 449572 48039
rect 453580 48078 453632 48084
rect 453946 48104 454002 48113
rect 452290 48039 452346 48048
rect 453946 48039 454002 48048
rect 450636 48010 450688 48016
rect 451280 47456 451332 47462
rect 450082 47424 450138 47433
rect 449532 47388 449584 47394
rect 450082 47359 450138 47368
rect 450450 47424 450506 47433
rect 450450 47359 450506 47368
rect 451278 47424 451280 47433
rect 451332 47424 451334 47433
rect 451334 47382 451412 47410
rect 451278 47359 451334 47368
rect 449532 47330 449584 47336
rect 447508 47252 447560 47258
rect 447508 47194 447560 47200
rect 446404 47048 446456 47054
rect 446404 46990 446456 46996
rect 446416 46510 446444 46990
rect 446404 46504 446456 46510
rect 446404 46446 446456 46452
rect 445300 46436 445352 46442
rect 445300 46378 445352 46384
rect 420000 45348 420052 45354
rect 420000 45290 420052 45296
rect 447520 45286 447548 47194
rect 449544 45490 449572 47330
rect 450096 45558 450124 47359
rect 450464 47326 450492 47359
rect 450452 47320 450504 47326
rect 450452 47262 450504 47268
rect 451280 47184 451332 47190
rect 451280 47126 451332 47132
rect 450084 45552 450136 45558
rect 450084 45494 450136 45500
rect 449532 45484 449584 45490
rect 449532 45426 449584 45432
rect 451292 45422 451320 47126
rect 451280 45416 451332 45422
rect 451280 45358 451332 45364
rect 451384 45354 451412 47382
rect 452304 47190 452332 48039
rect 452292 47184 452344 47190
rect 452292 47126 452344 47132
rect 453960 46986 453988 48039
rect 454604 47938 454632 48175
rect 455892 48006 455920 48175
rect 456996 48113 457024 49807
rect 458100 48210 458128 49807
rect 478564 49807 478566 49816
rect 480902 49872 480958 49881
rect 480902 49807 480958 49816
rect 478512 49778 478564 49784
rect 480916 49774 480944 49807
rect 480904 49768 480956 49774
rect 473358 49736 473414 49745
rect 480904 49710 480956 49716
rect 488262 49736 488318 49745
rect 473358 49671 473414 49680
rect 488262 49671 488318 49680
rect 495898 49736 495954 49745
rect 495898 49671 495900 49680
rect 459466 49056 459522 49065
rect 459466 48991 459522 49000
rect 459480 48278 459508 48991
rect 459928 48816 459980 48822
rect 459928 48758 459980 48764
rect 458364 48272 458416 48278
rect 458362 48240 458364 48249
rect 459468 48272 459520 48278
rect 458416 48240 458418 48249
rect 458088 48204 458140 48210
rect 459468 48214 459520 48220
rect 458362 48175 458418 48184
rect 458088 48146 458140 48152
rect 456982 48104 457038 48113
rect 456982 48039 457038 48048
rect 455880 48000 455932 48006
rect 455880 47942 455932 47948
rect 454592 47932 454644 47938
rect 454592 47874 454644 47880
rect 459940 47705 459968 48758
rect 461674 48240 461730 48249
rect 461674 48175 461730 48184
rect 462778 48240 462834 48249
rect 462778 48175 462834 48184
rect 463514 48240 463570 48249
rect 463514 48175 463570 48184
rect 463882 48240 463938 48249
rect 463882 48175 463938 48184
rect 465170 48240 465226 48249
rect 465170 48175 465226 48184
rect 465906 48240 465962 48249
rect 465906 48175 465962 48184
rect 466274 48240 466330 48249
rect 466274 48175 466330 48184
rect 467562 48240 467618 48249
rect 467562 48175 467618 48184
rect 468298 48240 468354 48249
rect 468298 48175 468354 48184
rect 468666 48240 468722 48249
rect 468666 48175 468722 48184
rect 469218 48240 469274 48249
rect 469218 48175 469274 48184
rect 470874 48240 470930 48249
rect 470874 48175 470930 48184
rect 471242 48240 471298 48249
rect 471242 48175 471298 48184
rect 472162 48240 472218 48249
rect 472162 48175 472218 48184
rect 461688 47734 461716 48175
rect 461676 47728 461728 47734
rect 459926 47696 459982 47705
rect 461676 47670 461728 47676
rect 462792 47666 462820 48175
rect 459926 47631 459982 47640
rect 462780 47660 462832 47666
rect 462780 47602 462832 47608
rect 453948 46980 454000 46986
rect 453948 46922 454000 46928
rect 453960 46578 453988 46922
rect 463528 46646 463556 48175
rect 463896 47122 463924 48175
rect 463884 47116 463936 47122
rect 463884 47058 463936 47064
rect 465184 47054 465212 48175
rect 465172 47048 465224 47054
rect 465172 46990 465224 46996
rect 465920 46714 465948 48175
rect 466288 47258 466316 48175
rect 467576 47394 467604 48175
rect 467564 47388 467616 47394
rect 467564 47330 467616 47336
rect 466276 47252 466328 47258
rect 466276 47194 466328 47200
rect 468312 46782 468340 48175
rect 468680 47326 468708 48175
rect 469128 48136 469180 48142
rect 469126 48104 469128 48113
rect 469180 48104 469182 48113
rect 469126 48039 469182 48048
rect 469232 47462 469260 48175
rect 469220 47456 469272 47462
rect 469220 47398 469272 47404
rect 468668 47320 468720 47326
rect 468668 47262 468720 47268
rect 470888 46850 470916 48175
rect 471256 47190 471284 48175
rect 471244 47184 471296 47190
rect 471244 47126 471296 47132
rect 472176 46986 472204 48175
rect 473372 47598 473400 49671
rect 488276 48890 488304 49671
rect 495952 49671 495954 49680
rect 503534 49736 503590 49745
rect 503534 49671 503590 49680
rect 495900 49642 495952 49648
rect 503548 49638 503576 49671
rect 503536 49632 503588 49638
rect 493414 49600 493470 49609
rect 493414 49535 493470 49544
rect 498474 49600 498530 49609
rect 498474 49535 498530 49544
rect 500958 49600 501014 49609
rect 503536 49574 503588 49580
rect 505926 49600 505982 49609
rect 500958 49535 500960 49544
rect 493428 48958 493456 49535
rect 498488 49502 498516 49535
rect 501012 49535 501014 49544
rect 505926 49535 505982 49544
rect 508502 49600 508558 49609
rect 508502 49535 508558 49544
rect 510986 49600 511042 49609
rect 510986 49535 511042 49544
rect 513378 49600 513434 49609
rect 513378 49535 513434 49544
rect 515862 49600 515918 49609
rect 515862 49535 515918 49544
rect 520922 49600 520978 49609
rect 520922 49535 520978 49544
rect 525890 49600 525946 49609
rect 525890 49535 525946 49544
rect 500960 49506 501012 49512
rect 498476 49496 498528 49502
rect 498476 49438 498528 49444
rect 505940 49434 505968 49535
rect 505928 49428 505980 49434
rect 505928 49370 505980 49376
rect 508516 49366 508544 49535
rect 508504 49360 508556 49366
rect 508504 49302 508556 49308
rect 511000 49298 511028 49535
rect 510988 49292 511040 49298
rect 510988 49234 511040 49240
rect 513392 49162 513420 49535
rect 515876 49230 515904 49535
rect 515864 49224 515916 49230
rect 515864 49166 515916 49172
rect 513380 49156 513432 49162
rect 513380 49098 513432 49104
rect 520936 49094 520964 49535
rect 520924 49088 520976 49094
rect 520924 49030 520976 49036
rect 525904 49026 525932 49535
rect 525892 49020 525944 49026
rect 525892 48962 525944 48968
rect 493416 48952 493468 48958
rect 493416 48894 493468 48900
rect 488264 48884 488316 48890
rect 488264 48826 488316 48832
rect 478052 48272 478104 48278
rect 474370 48240 474426 48249
rect 474370 48175 474426 48184
rect 475658 48240 475714 48249
rect 475658 48175 475714 48184
rect 476946 48240 477002 48249
rect 476946 48175 476948 48184
rect 474384 48006 474412 48175
rect 475672 48142 475700 48175
rect 477000 48175 477002 48184
rect 478050 48240 478052 48249
rect 478104 48240 478106 48249
rect 478050 48175 478106 48184
rect 476948 48146 477000 48152
rect 475660 48136 475712 48142
rect 475660 48078 475712 48084
rect 474372 48000 474424 48006
rect 474372 47942 474424 47948
rect 473360 47592 473412 47598
rect 473360 47534 473412 47540
rect 472164 46980 472216 46986
rect 472164 46922 472216 46928
rect 470876 46844 470928 46850
rect 470876 46786 470928 46792
rect 468300 46776 468352 46782
rect 468300 46718 468352 46724
rect 465908 46708 465960 46714
rect 465908 46650 465960 46656
rect 463516 46640 463568 46646
rect 463516 46582 463568 46588
rect 453948 46572 454000 46578
rect 453948 46514 454000 46520
rect 451372 45348 451424 45354
rect 451372 45290 451424 45296
rect 416504 45280 416556 45286
rect 416504 45222 416556 45228
rect 447508 45280 447560 45286
rect 447508 45222 447560 45228
rect 494704 44872 494756 44878
rect 494704 44814 494756 44820
rect 483664 43444 483716 43450
rect 483664 43386 483716 43392
rect 431960 37936 432012 37942
rect 431960 37878 432012 37884
rect 420920 35216 420972 35222
rect 420920 35158 420972 35164
rect 416780 17264 416832 17270
rect 416780 17206 416832 17212
rect 416792 16574 416820 17206
rect 407132 16546 407252 16574
rect 409892 16546 410840 16574
rect 414032 16546 414336 16574
rect 416792 16546 417464 16574
rect 403624 3936 403676 3942
rect 403624 3878 403676 3884
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 403636 480 403664 3878
rect 407224 480 407252 16546
rect 410812 480 410840 16546
rect 414308 480 414336 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 35158
rect 427820 22772 427872 22778
rect 427820 22714 427872 22720
rect 423680 21412 423732 21418
rect 423680 21354 423732 21360
rect 423692 2786 423720 21354
rect 427832 16574 427860 22714
rect 431972 16574 432000 37878
rect 473360 32428 473412 32434
rect 473360 32370 473412 32376
rect 445760 31068 445812 31074
rect 445760 31010 445812 31016
rect 441620 29640 441672 29646
rect 441620 29582 441672 29588
rect 434720 28280 434772 28286
rect 434720 28222 434772 28228
rect 434732 16574 434760 28222
rect 438860 25560 438912 25566
rect 438860 25502 438912 25508
rect 438872 16574 438900 25502
rect 441632 16574 441660 29582
rect 427832 16546 428504 16574
rect 431972 16546 432092 16574
rect 434732 16546 435128 16574
rect 438872 16546 439176 16574
rect 441632 16546 442672 16574
rect 423680 2780 423732 2786
rect 423680 2722 423732 2728
rect 424968 2780 425020 2786
rect 424968 2722 425020 2728
rect 424980 480 425008 2722
rect 428476 480 428504 16546
rect 432064 480 432092 16546
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 439148 480 439176 16546
rect 442644 480 442672 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 31010
rect 456800 26920 456852 26926
rect 456800 26862 456852 26868
rect 448520 24132 448572 24138
rect 448520 24074 448572 24080
rect 448532 2786 448560 24074
rect 456812 16574 456840 26862
rect 473372 16574 473400 32370
rect 456812 16546 456932 16574
rect 473372 16546 474136 16574
rect 453304 3868 453356 3874
rect 453304 3810 453356 3816
rect 448520 2780 448572 2786
rect 448520 2722 448572 2728
rect 449808 2780 449860 2786
rect 449808 2722 449860 2728
rect 449820 480 449848 2722
rect 453316 480 453344 3810
rect 456904 480 456932 16546
rect 460388 3800 460440 3806
rect 460388 3742 460440 3748
rect 460400 480 460428 3742
rect 463976 3732 464028 3738
rect 463976 3674 464028 3680
rect 463988 480 464016 3674
rect 467472 3664 467524 3670
rect 467472 3606 467524 3612
rect 467484 480 467512 3606
rect 471060 3596 471112 3602
rect 471060 3538 471112 3544
rect 471072 480 471100 3538
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 481732 7608 481784 7614
rect 481732 7550 481784 7556
rect 478144 3528 478196 3534
rect 478144 3470 478196 3476
rect 478156 480 478184 3470
rect 481744 480 481772 7550
rect 483676 2922 483704 43386
rect 492312 10328 492364 10334
rect 492312 10270 492364 10276
rect 488816 8968 488868 8974
rect 488816 8910 488868 8916
rect 483664 2916 483716 2922
rect 483664 2858 483716 2864
rect 485228 2916 485280 2922
rect 485228 2858 485280 2864
rect 485240 480 485268 2858
rect 488828 480 488856 8910
rect 492324 480 492352 10270
rect 494716 3534 494744 44814
rect 512644 42084 512696 42090
rect 512644 42026 512696 42032
rect 502340 39364 502392 39370
rect 502340 39306 502392 39312
rect 502352 16574 502380 39306
rect 502352 16546 503024 16574
rect 498936 11756 498988 11762
rect 498936 11698 498988 11704
rect 494704 3528 494756 3534
rect 494704 3470 494756 3476
rect 495900 3528 495952 3534
rect 495900 3470 495952 3476
rect 495912 480 495940 3470
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 11698
rect 502996 480 503024 16546
rect 506480 14476 506532 14482
rect 506480 14418 506532 14424
rect 506492 480 506520 14418
rect 508504 13116 508556 13122
rect 508504 13058 508556 13064
rect 508516 4146 508544 13058
rect 508504 4140 508556 4146
rect 508504 4082 508556 4088
rect 510068 4140 510120 4146
rect 510068 4082 510120 4088
rect 510080 480 510108 4082
rect 512656 3534 512684 42026
rect 523040 40724 523092 40730
rect 523040 40666 523092 40672
rect 523052 16574 523080 40666
rect 547880 36576 547932 36582
rect 547880 36518 547932 36524
rect 547892 16574 547920 36518
rect 555424 33788 555476 33794
rect 555424 33730 555476 33736
rect 523052 16546 523816 16574
rect 547892 16546 548656 16574
rect 517152 5296 517204 5302
rect 517152 5238 517204 5244
rect 512644 3528 512696 3534
rect 512644 3470 512696 3476
rect 513564 3528 513616 3534
rect 513564 3470 513616 3476
rect 513576 480 513604 3470
rect 517164 480 517192 5238
rect 520740 5228 520792 5234
rect 520740 5170 520792 5176
rect 520752 480 520780 5170
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 527824 5160 527876 5166
rect 527824 5102 527876 5108
rect 527836 480 527864 5102
rect 531320 5092 531372 5098
rect 531320 5034 531372 5040
rect 531332 480 531360 5034
rect 534908 5024 534960 5030
rect 534908 4966 534960 4972
rect 534920 480 534948 4966
rect 538404 4956 538456 4962
rect 538404 4898 538456 4904
rect 538416 480 538444 4898
rect 541992 4888 542044 4894
rect 541992 4830 542044 4836
rect 542004 480 542032 4830
rect 545488 4820 545540 4826
rect 545488 4762 545540 4768
rect 545500 480 545528 4762
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 552664 6316 552716 6322
rect 552664 6258 552716 6264
rect 552676 480 552704 6258
rect 555436 3534 555464 33730
rect 555424 3528 555476 3534
rect 555424 3470 555476 3476
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556172 480 556200 3470
rect 558196 2922 558224 246366
rect 558932 240802 558960 329151
rect 563716 325650 563744 461042
rect 576124 461032 576176 461038
rect 576124 460974 576176 460980
rect 563794 459640 563850 459649
rect 563794 459575 563850 459584
rect 563808 405686 563836 459575
rect 563796 405680 563848 405686
rect 563796 405622 563848 405628
rect 576136 379506 576164 460974
rect 576124 379500 576176 379506
rect 576124 379442 576176 379448
rect 563704 325644 563756 325650
rect 563704 325586 563756 325592
rect 576124 246356 576176 246362
rect 576124 246298 576176 246304
rect 558840 240786 558960 240802
rect 558828 240780 558960 240786
rect 558880 240774 558960 240780
rect 558828 240722 558880 240728
rect 562324 238128 562376 238134
rect 562324 238070 562376 238076
rect 558918 229256 558974 229265
rect 558918 229191 558974 229200
rect 558932 129713 558960 229191
rect 558918 129704 558974 129713
rect 558918 129639 558974 129648
rect 559564 110424 559616 110430
rect 559564 110366 559616 110372
rect 559576 99006 559604 110366
rect 559564 99000 559616 99006
rect 559564 98942 559616 98948
rect 562336 2922 562364 238070
rect 565084 99000 565136 99006
rect 565084 98942 565136 98948
rect 565096 91798 565124 98942
rect 565084 91792 565136 91798
rect 565084 91734 565136 91740
rect 569960 91792 570012 91798
rect 569960 91734 570012 91740
rect 569972 85542 570000 91734
rect 569960 85536 570012 85542
rect 569960 85478 570012 85484
rect 573364 85536 573416 85542
rect 573364 85478 573416 85484
rect 573376 73166 573404 85478
rect 573364 73160 573416 73166
rect 573364 73102 573416 73108
rect 563060 15904 563112 15910
rect 563060 15846 563112 15852
rect 558184 2916 558236 2922
rect 558184 2858 558236 2864
rect 559748 2916 559800 2922
rect 559748 2858 559800 2864
rect 562324 2916 562376 2922
rect 562324 2858 562376 2864
rect 559760 480 559788 2858
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 15846
rect 570328 6248 570380 6254
rect 570328 6190 570380 6196
rect 566832 2916 566884 2922
rect 566832 2858 566884 2864
rect 566844 480 566872 2858
rect 570340 480 570368 6190
rect 573916 6180 573968 6186
rect 573916 6122 573968 6128
rect 573928 480 573956 6122
rect 576136 4146 576164 246298
rect 577516 100706 577544 466482
rect 577596 465180 577648 465186
rect 577596 465122 577648 465128
rect 577608 139398 577636 465122
rect 577700 179382 577728 466822
rect 577872 466812 577924 466818
rect 577872 466754 577924 466760
rect 577780 466608 577832 466614
rect 577780 466550 577832 466556
rect 577792 193186 577820 466550
rect 577884 219230 577912 466754
rect 577964 466744 578016 466750
rect 577964 466686 578016 466692
rect 577976 233238 578004 466686
rect 580540 466676 580592 466682
rect 580540 466618 580592 466624
rect 580264 466472 580316 466478
rect 580264 466414 580316 466420
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 579986 454472 580042 454481
rect 579986 454407 580042 454416
rect 579620 325644 579672 325650
rect 579620 325586 579672 325592
rect 579632 325281 579660 325586
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 580000 312089 580028 454407
rect 580170 454336 580226 454345
rect 580170 454271 580226 454280
rect 580080 431928 580132 431934
rect 580080 431870 580132 431876
rect 580092 431633 580120 431870
rect 580078 431624 580134 431633
rect 580078 431559 580134 431568
rect 580080 419484 580132 419490
rect 580080 419426 580132 419432
rect 580092 418305 580120 419426
rect 580078 418296 580134 418305
rect 580078 418231 580134 418240
rect 580080 405680 580132 405686
rect 580080 405622 580132 405628
rect 580092 404977 580120 405622
rect 580078 404968 580134 404977
rect 580078 404903 580134 404912
rect 580080 379500 580132 379506
rect 580080 379442 580132 379448
rect 580092 378457 580120 379442
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580080 353252 580132 353258
rect 580080 353194 580132 353200
rect 580092 351937 580120 353194
rect 580078 351928 580134 351937
rect 580078 351863 580134 351872
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580184 298761 580212 454271
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 578884 233912 578936 233918
rect 578884 233854 578936 233860
rect 577964 233232 578016 233238
rect 577964 233174 578016 233180
rect 577872 219224 577924 219230
rect 577872 219166 577924 219172
rect 577780 193180 577832 193186
rect 577780 193122 577832 193128
rect 577688 179376 577740 179382
rect 577688 179318 577740 179324
rect 577596 139392 577648 139398
rect 577596 139334 577648 139340
rect 577504 100700 577556 100706
rect 577504 100642 577556 100648
rect 576124 4140 576176 4146
rect 576124 4082 576176 4088
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 578896 3262 578924 233854
rect 579620 233232 579672 233238
rect 579620 233174 579672 233180
rect 579632 232393 579660 233174
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579988 219224 580040 219230
rect 579988 219166 580040 219172
rect 580000 219065 580028 219166
rect 579986 219056 580042 219065
rect 579986 218991 580042 219000
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 580080 179376 580132 179382
rect 580080 179318 580132 179324
rect 580092 179217 580120 179318
rect 580078 179208 580134 179217
rect 580078 179143 580134 179152
rect 579620 139392 579672 139398
rect 579618 139360 579620 139369
rect 579672 139360 579674 139369
rect 579618 139295 579674 139304
rect 580276 112849 580304 466414
rect 580356 465112 580408 465118
rect 580356 465054 580408 465060
rect 580368 152697 580396 465054
rect 580448 463752 580500 463758
rect 580448 463694 580500 463700
rect 580460 205737 580488 463694
rect 580552 245585 580580 466618
rect 580724 460964 580776 460970
rect 580724 460906 580776 460912
rect 580630 454200 580686 454209
rect 580630 454135 580686 454144
rect 580644 258913 580672 454135
rect 580736 365129 580764 460906
rect 580814 454880 580870 454889
rect 580814 454815 580870 454824
rect 580722 365120 580778 365129
rect 580722 365055 580778 365064
rect 580828 272241 580856 454815
rect 580814 272232 580870 272241
rect 580814 272167 580870 272176
rect 580630 258904 580686 258913
rect 580630 258839 580686 258848
rect 580538 245576 580594 245585
rect 580538 245511 580594 245520
rect 580540 238060 580592 238066
rect 580540 238002 580592 238008
rect 580446 205728 580502 205737
rect 580446 205663 580502 205672
rect 580552 165889 580580 238002
rect 582380 236700 582432 236706
rect 582380 236642 582432 236648
rect 580538 165880 580594 165889
rect 580538 165815 580594 165824
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 580448 134700 580500 134706
rect 580448 134642 580500 134648
rect 580356 134564 580408 134570
rect 580356 134506 580408 134512
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 579712 100700 579764 100706
rect 579712 100642 579764 100648
rect 579724 99521 579752 100642
rect 579710 99512 579766 99521
rect 579710 99447 579766 99456
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580368 59673 580396 134506
rect 580460 86193 580488 134642
rect 580908 134632 580960 134638
rect 580908 134574 580960 134580
rect 580920 126041 580948 134574
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 580446 86184 580502 86193
rect 580446 86119 580502 86128
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 582392 16574 582420 236642
rect 582392 16546 583432 16574
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 578884 3256 578936 3262
rect 578884 3198 578936 3204
rect 581012 480 581040 3402
rect 582196 3256 582248 3262
rect 582196 3198 582248 3204
rect 582208 480 582236 3198
rect 583404 480 583432 16546
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3330 501744 3386 501800
rect 3514 514800 3570 514856
rect 3422 475632 3478 475688
rect 30102 680312 30158 680368
rect 34886 680448 34942 680504
rect 46846 682624 46902 682680
rect 53654 682352 53710 682408
rect 51630 682216 51686 682272
rect 60738 680992 60794 681048
rect 75550 681944 75606 682000
rect 137742 682080 137798 682136
rect 168838 681808 168894 681864
rect 169758 679768 169814 679824
rect 197174 682488 197230 682544
rect 195150 682080 195206 682136
rect 192758 681944 192814 682000
rect 144274 679632 144330 679688
rect 79046 679496 79102 679552
rect 190044 679224 190100 679280
rect 3238 462576 3294 462632
rect 3238 423544 3294 423600
rect 3330 410488 3386 410544
rect 3606 452784 3662 452840
rect 3514 449540 3570 449576
rect 3514 449520 3516 449540
rect 3516 449520 3568 449540
rect 3568 449520 3570 449540
rect 3514 449384 3570 449440
rect 3422 358400 3478 358456
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 4066 397432 4122 397488
rect 3974 371320 4030 371376
rect 3882 319232 3938 319288
rect 3790 306176 3846 306232
rect 3698 293120 3754 293176
rect 3606 267144 3662 267200
rect 3514 254088 3570 254144
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3422 58520 3478 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 14738 449928 14794 449984
rect 15106 451968 15162 452024
rect 17222 385872 17278 385928
rect 16762 380976 16818 381032
rect 16946 359896 17002 359952
rect 16854 283736 16910 283792
rect 16762 281016 16818 281072
rect 16762 186904 16818 186960
rect 17038 358264 17094 358320
rect 16946 260752 17002 260808
rect 17130 285776 17186 285832
rect 16854 183776 16910 183832
rect 16762 86808 16818 86864
rect 17590 386824 17646 386880
rect 17314 379888 17370 379944
rect 17222 285640 17278 285696
rect 17406 378120 17462 378176
rect 17314 279928 17370 279984
rect 17590 286864 17646 286920
rect 17590 285776 17646 285832
rect 17498 283736 17554 283792
rect 17590 282784 17646 282840
rect 17774 378120 17830 378176
rect 17774 285640 17830 285696
rect 17498 281016 17554 281072
rect 17406 278704 17462 278760
rect 17130 186904 17186 186960
rect 17130 185952 17186 186008
rect 16946 83680 17002 83736
rect 17406 260752 17462 260808
rect 17406 259936 17462 259992
rect 17314 258304 17370 258360
rect 17222 179424 17278 179480
rect 17682 278704 17738 278760
rect 17682 278160 17738 278216
rect 17590 182824 17646 182880
rect 17498 181056 17554 181112
rect 17406 159976 17462 160032
rect 17314 158344 17370 158400
rect 17130 85856 17186 85912
rect 18786 385872 18842 385928
rect 18878 383696 18934 383752
rect 18970 382744 19026 382800
rect 19062 380976 19118 381032
rect 19154 359896 19210 359952
rect 134338 449656 134394 449712
rect 151082 435240 151138 435296
rect 156602 450064 156658 450120
rect 19338 386824 19394 386880
rect 19246 357992 19302 358048
rect 91006 349832 91062 349888
rect 93490 349832 93546 349888
rect 98550 349832 98606 349888
rect 103518 349832 103574 349888
rect 38474 349560 38530 349616
rect 50802 349560 50858 349616
rect 56046 349560 56102 349616
rect 58530 349560 58586 349616
rect 61106 349560 61162 349616
rect 62854 349560 62910 349616
rect 68742 349560 68798 349616
rect 72238 349560 72294 349616
rect 53654 349016 53710 349072
rect 17866 258168 17922 258224
rect 18694 249736 18750 249792
rect 17774 185952 17830 186008
rect 17866 179968 17922 180024
rect 17866 179424 17922 179480
rect 17774 178200 17830 178256
rect 17590 82864 17646 82920
rect 17498 80960 17554 81016
rect 17866 79872 17922 79928
rect 17774 78104 17830 78160
rect 17406 59880 17462 59936
rect 17314 58248 17370 58304
rect 62026 349052 62028 349072
rect 62028 349052 62080 349072
rect 62080 349052 62082 349072
rect 62026 349016 62082 349052
rect 36174 347656 36230 347712
rect 39578 347656 39634 347712
rect 42798 347692 42800 347712
rect 42800 347692 42852 347712
rect 42852 347692 42854 347712
rect 42798 347656 42854 347692
rect 44178 347656 44234 347712
rect 45374 347656 45430 347712
rect 18786 146784 18842 146840
rect 18786 47912 18842 47968
rect 18694 47776 18750 47832
rect 19614 247968 19670 248024
rect 19430 147328 19486 147384
rect 37186 347248 37242 347304
rect 46570 347676 46626 347712
rect 46570 347656 46572 347676
rect 46572 347656 46624 347676
rect 46624 347656 46626 347676
rect 47582 347656 47638 347712
rect 48594 347656 48650 347712
rect 50066 347656 50122 347712
rect 51262 347656 51318 347712
rect 52366 347656 52422 347712
rect 53470 347656 53526 347712
rect 41786 346840 41842 346896
rect 41326 346432 41382 346488
rect 63682 347656 63738 347712
rect 64786 347692 64788 347712
rect 64788 347692 64840 347712
rect 64840 347692 64842 347712
rect 64786 347656 64842 347692
rect 65154 347676 65210 347712
rect 65154 347656 65156 347676
rect 65156 347656 65208 347676
rect 65208 347656 65210 347676
rect 56598 347384 56654 347440
rect 59358 347384 59414 347440
rect 60830 347384 60886 347440
rect 55126 346704 55182 346760
rect 41786 345208 41842 345264
rect 42706 345208 42762 345264
rect 57978 347112 58034 347168
rect 60738 347112 60794 347168
rect 57978 346432 58034 346488
rect 61934 347112 61990 347168
rect 65982 347656 66038 347712
rect 66258 347676 66314 347712
rect 66258 347656 66260 347676
rect 66260 347656 66312 347676
rect 66312 347656 66314 347676
rect 68374 349016 68430 349072
rect 67730 347656 67786 347712
rect 71134 347656 71190 347712
rect 74354 348472 74410 348528
rect 78494 349016 78550 349072
rect 86038 349016 86094 349072
rect 73250 347656 73306 347712
rect 73710 347656 73766 347712
rect 75458 347656 75514 347712
rect 76102 347656 76158 347712
rect 76746 347656 76802 347712
rect 78034 347656 78090 347712
rect 79138 347656 79194 347712
rect 81070 347656 81126 347712
rect 83646 347656 83702 347712
rect 96066 347656 96122 347712
rect 100942 347656 100998 347712
rect 106094 347656 106150 347712
rect 108670 347656 108726 347712
rect 111062 347656 111118 347712
rect 113454 347656 113510 347712
rect 115846 347656 115902 347712
rect 118606 347656 118662 347712
rect 120998 347656 121054 347712
rect 123390 347656 123446 347712
rect 125966 347656 126022 347712
rect 69294 347112 69350 347168
rect 75458 346432 75514 346488
rect 150990 335416 151046 335472
rect 93490 249736 93546 249792
rect 95882 249736 95938 249792
rect 98550 249736 98606 249792
rect 103518 249736 103574 249792
rect 106002 249736 106058 249792
rect 108578 249736 108634 249792
rect 111062 249756 111118 249792
rect 111062 249736 111064 249756
rect 111064 249736 111116 249756
rect 111116 249736 111118 249756
rect 50802 249600 50858 249656
rect 53654 249600 53710 249656
rect 56046 249600 56102 249656
rect 58530 249600 58586 249656
rect 113454 249600 113510 249656
rect 115846 249600 115902 249656
rect 120906 249600 120962 249656
rect 35898 248240 35954 248296
rect 36450 248276 36452 248296
rect 36452 248276 36504 248296
rect 36504 248276 36506 248296
rect 36450 248240 36506 248276
rect 38658 248260 38714 248296
rect 38658 248240 38660 248260
rect 38660 248240 38712 248260
rect 38712 248240 38714 248260
rect 44178 248240 44234 248296
rect 46662 248260 46718 248296
rect 46662 248240 46664 248260
rect 46664 248240 46716 248260
rect 46716 248240 46718 248260
rect 50158 248240 50214 248296
rect 61198 248240 61254 248296
rect 61382 248240 61438 248296
rect 62118 248240 62174 248296
rect 63590 248276 63592 248296
rect 63592 248276 63644 248296
rect 63644 248276 63646 248296
rect 63590 248240 63646 248276
rect 64878 248260 64934 248296
rect 64878 248240 64880 248260
rect 64880 248240 64932 248260
rect 64932 248240 64934 248260
rect 37278 248124 37334 248160
rect 37278 248104 37280 248124
rect 37280 248104 37332 248124
rect 37332 248104 37334 248124
rect 40038 248104 40094 248160
rect 41418 248124 41474 248160
rect 41418 248104 41420 248124
rect 41420 248104 41472 248124
rect 41472 248104 41474 248124
rect 29550 247696 29606 247752
rect 43074 248104 43130 248160
rect 45282 248104 45338 248160
rect 47582 248104 47638 248160
rect 48686 247832 48742 247888
rect 65982 248240 66038 248296
rect 67638 248240 67694 248296
rect 70950 248240 71006 248296
rect 73802 248260 73858 248296
rect 73802 248240 73804 248260
rect 73804 248240 73856 248260
rect 73856 248240 73858 248260
rect 63498 247988 63554 248024
rect 63498 247968 63500 247988
rect 63500 247968 63552 247988
rect 63552 247968 63554 247988
rect 58070 247832 58126 247888
rect 59450 247832 59506 247888
rect 66258 247852 66314 247888
rect 77298 248240 77354 248296
rect 78494 248240 78550 248296
rect 83646 248240 83702 248296
rect 81070 247968 81126 248024
rect 66258 247832 66260 247852
rect 66260 247832 66312 247852
rect 66312 247832 66314 247852
rect 38106 247560 38162 247616
rect 52366 247424 52422 247480
rect 67730 247832 67786 247888
rect 68374 247832 68430 247888
rect 76102 247832 76158 247888
rect 74998 247696 75054 247752
rect 75918 247716 75974 247752
rect 75918 247696 75920 247716
rect 75920 247696 75972 247716
rect 75972 247696 75974 247716
rect 52366 247016 52422 247072
rect 53746 247288 53802 247344
rect 55126 247016 55182 247072
rect 56506 247016 56562 247072
rect 71778 247560 71834 247616
rect 86038 247968 86094 248024
rect 88246 247968 88302 248024
rect 91006 247968 91062 248024
rect 101218 247968 101274 248024
rect 69018 247424 69074 247480
rect 70398 247308 70454 247344
rect 70398 247288 70400 247308
rect 70400 247288 70452 247308
rect 70452 247288 70454 247308
rect 73250 247288 73306 247344
rect 73158 247172 73214 247208
rect 73158 247152 73160 247172
rect 73160 247152 73212 247172
rect 73212 247152 73214 247172
rect 57978 247016 58034 247072
rect 63222 247016 63278 247072
rect 150438 234660 150494 234696
rect 150438 234640 150440 234660
rect 150440 234640 150492 234660
rect 150492 234640 150494 234660
rect 48318 149504 48374 149560
rect 50802 149504 50858 149560
rect 56046 149504 56102 149560
rect 58530 149504 58586 149560
rect 60646 149504 60702 149560
rect 71226 149504 71282 149560
rect 73618 149504 73674 149560
rect 83554 149504 83610 149560
rect 93490 149504 93546 149560
rect 98550 149504 98606 149560
rect 103518 149504 103574 149560
rect 113454 149504 113510 149560
rect 115846 149504 115902 149560
rect 120906 149504 120962 149560
rect 53654 148960 53710 149016
rect 19522 147192 19578 147248
rect 19522 48048 19578 48104
rect 18970 47504 19026 47560
rect 35898 147600 35954 147656
rect 37002 147620 37058 147656
rect 37002 147600 37004 147620
rect 37004 147600 37056 147620
rect 37056 147600 37058 147620
rect 38106 147600 38162 147656
rect 39578 147600 39634 147656
rect 43074 147600 43130 147656
rect 44178 147600 44234 147656
rect 45282 147600 45338 147656
rect 46570 147600 46626 147656
rect 47674 147600 47730 147656
rect 48686 147600 48742 147656
rect 50158 147620 50214 147656
rect 50158 147600 50160 147620
rect 50160 147600 50212 147620
rect 50212 147600 50214 147620
rect 51446 147600 51502 147656
rect 52274 147600 52330 147656
rect 53378 147600 53434 147656
rect 54022 147600 54078 147656
rect 56046 147600 56102 147656
rect 58070 147600 58126 147656
rect 59542 147636 59544 147656
rect 59544 147636 59596 147656
rect 59596 147636 59598 147656
rect 59542 147600 59598 147636
rect 61658 147600 61714 147656
rect 62762 147600 62818 147656
rect 63590 147620 63646 147656
rect 63590 147600 63592 147620
rect 63592 147600 63644 147620
rect 63644 147600 63646 147620
rect 60646 147464 60702 147520
rect 63866 147600 63922 147656
rect 65154 147600 65210 147656
rect 66166 147600 66222 147656
rect 66350 147600 66406 147656
rect 67638 147600 67694 147656
rect 68282 147600 68338 147656
rect 68466 147600 68522 147656
rect 69754 147600 69810 147656
rect 70398 147192 70454 147248
rect 71042 147192 71098 147248
rect 76102 148960 76158 149016
rect 86038 148960 86094 149016
rect 72146 147600 72202 147656
rect 73250 147600 73306 147656
rect 73710 147600 73766 147656
rect 75642 147600 75698 147656
rect 76930 147600 76986 147656
rect 78034 147600 78090 147656
rect 78494 147600 78550 147656
rect 79138 147600 79194 147656
rect 81070 147600 81126 147656
rect 88246 147600 88302 147656
rect 91006 147600 91062 147656
rect 95974 147600 96030 147656
rect 100942 147600 100998 147656
rect 75826 147464 75882 147520
rect 106094 147600 106150 147656
rect 108854 147600 108910 147656
rect 111614 147600 111670 147656
rect 157982 456320 158038 456376
rect 157890 452240 157946 452296
rect 156786 450472 156842 450528
rect 156786 147464 156842 147520
rect 158166 455504 158222 455560
rect 158534 451560 158590 451616
rect 158810 429256 158866 429312
rect 158810 329704 158866 329760
rect 158718 229200 158774 229256
rect 151266 135768 151322 135824
rect 158718 129648 158774 129704
rect 53470 49852 53472 49872
rect 53472 49852 53524 49872
rect 53524 49852 53526 49872
rect 53470 49816 53526 49852
rect 48318 49544 48374 49600
rect 50802 49544 50858 49600
rect 36818 48220 36820 48240
rect 36820 48220 36872 48240
rect 36872 48220 36874 48240
rect 36818 48184 36874 48220
rect 43166 48184 43222 48240
rect 44178 48184 44234 48240
rect 45374 48184 45430 48240
rect 46570 48184 46626 48240
rect 47582 48184 47638 48240
rect 48686 48184 48742 48240
rect 49698 48184 49754 48240
rect 50250 48184 50306 48240
rect 51446 48184 51502 48240
rect 52366 48184 52422 48240
rect 60646 49816 60702 49872
rect 53654 49544 53710 49600
rect 56046 49544 56102 49600
rect 58530 49544 58586 49600
rect 54574 48184 54630 48240
rect 55862 48184 55918 48240
rect 57978 48184 58034 48240
rect 59542 48220 59544 48240
rect 59544 48220 59596 48240
rect 59596 48220 59598 48240
rect 59542 48184 59598 48220
rect 57058 47504 57114 47560
rect 91006 49680 91062 49736
rect 95882 49700 95938 49736
rect 95882 49680 95884 49700
rect 95884 49680 95936 49700
rect 95936 49680 95938 49700
rect 80978 49544 81034 49600
rect 83554 49544 83610 49600
rect 86038 49544 86094 49600
rect 88246 49564 88302 49600
rect 88246 49544 88248 49564
rect 88248 49544 88300 49564
rect 88300 49544 88302 49564
rect 98550 49544 98606 49600
rect 103518 49544 103574 49600
rect 106002 49544 106058 49600
rect 61198 48204 61254 48240
rect 61198 48184 61200 48204
rect 61200 48184 61252 48204
rect 61252 48184 61254 48204
rect 61382 48184 61438 48240
rect 62210 48184 62266 48240
rect 63958 48184 64014 48240
rect 65062 48184 65118 48240
rect 65982 48184 66038 48240
rect 66258 48184 66314 48240
rect 67638 48184 67694 48240
rect 68374 48184 68430 48240
rect 68558 48184 68614 48240
rect 69754 48184 69810 48240
rect 71134 48184 71190 48240
rect 71778 48184 71834 48240
rect 73250 48184 73306 48240
rect 73802 48184 73858 48240
rect 74354 48184 74410 48240
rect 76102 48184 76158 48240
rect 76378 48184 76434 48240
rect 78034 48220 78036 48240
rect 78036 48220 78088 48240
rect 78088 48220 78090 48240
rect 78034 48184 78090 48220
rect 78494 48184 78550 48240
rect 93582 48184 93638 48240
rect 100942 48184 100998 48240
rect 108854 48184 108910 48240
rect 111154 48184 111210 48240
rect 115846 48184 115902 48240
rect 118606 48184 118662 48240
rect 125966 48220 125968 48240
rect 125968 48220 126020 48240
rect 126020 48220 126022 48240
rect 125966 48184 126022 48220
rect 60646 47912 60702 47968
rect 63866 48048 63922 48104
rect 71042 48048 71098 48104
rect 163594 463936 163650 463992
rect 161018 49408 161074 49464
rect 163502 462304 163558 462360
rect 163962 463800 164018 463856
rect 163778 463664 163834 463720
rect 163870 456048 163926 456104
rect 166630 464072 166686 464128
rect 168010 454688 168066 454744
rect 170402 461488 170458 461544
rect 169114 460128 169170 460184
rect 169206 458768 169262 458824
rect 169574 452920 169630 452976
rect 174450 459856 174506 459912
rect 175186 459992 175242 460048
rect 175002 459720 175058 459776
rect 175094 349016 175150 349072
rect 174542 247968 174598 248024
rect 171782 247832 171838 247888
rect 183006 461352 183062 461408
rect 182822 461216 182878 461272
rect 180062 457680 180118 457736
rect 177762 448704 177818 448760
rect 180706 451696 180762 451752
rect 180706 248104 180762 248160
rect 182914 457136 182970 457192
rect 180154 147328 180210 147384
rect 183190 461080 183246 461136
rect 183098 459176 183154 459232
rect 183374 460944 183430 461000
rect 183190 148960 183246 149016
rect 185582 458632 185638 458688
rect 183466 450200 183522 450256
rect 183374 148824 183430 148880
rect 185766 459040 185822 459096
rect 185950 458496 186006 458552
rect 185858 454008 185914 454064
rect 187514 452104 187570 452160
rect 187422 449520 187478 449576
rect 188434 457000 188490 457056
rect 188710 456864 188766 456920
rect 189722 453192 189778 453248
rect 190274 452376 190330 452432
rect 190182 450608 190238 450664
rect 190366 451424 190422 451480
rect 190826 348608 190882 348664
rect 191102 450880 191158 450936
rect 190642 347384 190698 347440
rect 190642 347112 190698 347168
rect 190826 347540 190882 347576
rect 190826 347520 190828 347540
rect 190828 347520 190880 347540
rect 190880 347520 190882 347540
rect 191286 347520 191342 347576
rect 190826 347384 190882 347440
rect 195150 452648 195206 452704
rect 193218 451832 193274 451888
rect 191746 348608 191802 348664
rect 191654 347656 191710 347712
rect 191562 347384 191618 347440
rect 191470 347248 191526 347304
rect 193678 451424 193734 451480
rect 194782 452376 194838 452432
rect 194138 450336 194194 450392
rect 195886 452104 195942 452160
rect 197818 450608 197874 450664
rect 200670 454824 200726 454880
rect 201406 454280 201462 454336
rect 201038 454144 201094 454200
rect 202510 456184 202566 456240
rect 202142 454416 202198 454472
rect 203338 459584 203394 459640
rect 210422 450472 210478 450528
rect 231858 466520 231914 466576
rect 229006 452784 229062 452840
rect 227902 451832 227958 451888
rect 230110 451968 230166 452024
rect 232318 449928 232374 449984
rect 233882 454688 233938 454744
rect 234802 461488 234858 461544
rect 236090 680992 236146 681048
rect 237470 680312 237526 680368
rect 237562 679496 237618 679552
rect 240230 680448 240286 680504
rect 244462 682624 244518 682680
rect 247314 682352 247370 682408
rect 247130 682216 247186 682272
rect 250074 679768 250130 679824
rect 251546 462848 251602 462904
rect 229742 449792 229798 449848
rect 254122 678136 254178 678192
rect 255502 679632 255558 679688
rect 255594 457408 255650 457464
rect 280250 458904 280306 458960
rect 279054 449928 279110 449984
rect 280158 451696 280214 451752
rect 283010 455640 283066 455696
rect 283194 454552 283250 454608
rect 288714 462576 288770 462632
rect 284298 462440 284354 462496
rect 283930 454008 283986 454064
rect 285862 456048 285918 456104
rect 287610 457272 287666 457328
rect 289266 457136 289322 457192
rect 292026 457408 292082 457464
rect 291934 453464 291990 453520
rect 390650 682488 390706 682544
rect 390558 681944 390614 682000
rect 389178 678952 389234 679008
rect 296718 457136 296774 457192
rect 295246 451968 295302 452024
rect 300490 457544 300546 457600
rect 300398 453328 300454 453384
rect 302422 462712 302478 462768
rect 304814 455640 304870 455696
rect 303342 451560 303398 451616
rect 304446 453328 304502 453384
rect 305550 453192 305606 453248
rect 308494 451560 308550 451616
rect 309414 457680 309470 457736
rect 313646 452920 313702 452976
rect 315578 456048 315634 456104
rect 315118 452240 315174 452296
rect 318430 453056 318486 453112
rect 321098 460128 321154 460184
rect 322846 450472 322902 450528
rect 324502 458768 324558 458824
rect 327170 458768 327226 458824
rect 324318 452648 324374 452704
rect 326250 457000 326306 457056
rect 327630 453056 327686 453112
rect 330942 453192 330998 453248
rect 333610 458360 333666 458416
rect 332874 456864 332930 456920
rect 349158 464072 349214 464128
rect 342534 458632 342590 458688
rect 345386 458496 345442 458552
rect 344926 450744 344982 450800
rect 348330 459040 348386 459096
rect 354678 463936 354734 463992
rect 350814 450608 350870 450664
rect 352286 451832 352342 451888
rect 351550 450200 351606 450256
rect 353758 450336 353814 450392
rect 358818 463800 358874 463856
rect 357346 450880 357402 450936
rect 357898 456864 357954 456920
rect 358726 450200 358782 450256
rect 361578 463664 361634 463720
rect 360290 459992 360346 460048
rect 360014 451424 360070 451480
rect 360198 450064 360254 450120
rect 360842 455912 360898 455968
rect 364338 462304 364394 462360
rect 371238 461352 371294 461408
rect 363786 455776 363842 455832
rect 363234 455504 363290 455560
rect 366362 459856 366418 459912
rect 365994 456320 366050 456376
rect 366730 458224 366786 458280
rect 368938 459176 368994 459232
rect 372250 459720 372306 459776
rect 377034 461216 377090 461272
rect 375838 451696 375894 451752
rect 380990 461080 381046 461136
rect 383658 460944 383714 461000
rect 379518 455504 379574 455560
rect 378782 450064 378838 450120
rect 380254 452784 380310 452840
rect 382186 452920 382242 452976
rect 383474 454008 383530 454064
rect 383566 452104 383622 452160
rect 383474 451832 383530 451888
rect 384670 451832 384726 451888
rect 355598 449792 355654 449848
rect 386142 449656 386198 449712
rect 388442 450744 388498 450800
rect 386418 449692 386420 449712
rect 386420 449692 386472 449712
rect 386472 449692 386474 449712
rect 386418 449656 386474 449692
rect 193218 449520 193274 449576
rect 193954 449520 194010 449576
rect 387614 449520 387670 449576
rect 194046 449248 194102 449304
rect 191838 345072 191894 345128
rect 308586 250416 308642 250472
rect 388626 450608 388682 450664
rect 388534 347520 388590 347576
rect 388442 147328 388498 147384
rect 389270 455504 389326 455560
rect 388626 146512 388682 146568
rect 389362 248240 389418 248296
rect 390006 449520 390062 449576
rect 390006 359352 390062 359408
rect 390742 682080 390798 682136
rect 416778 536852 416834 536888
rect 416778 536832 416780 536852
rect 416780 536832 416832 536852
rect 416832 536832 416834 536852
rect 392674 453328 392730 453384
rect 392582 450336 392638 450392
rect 393962 453464 394018 453520
rect 392582 147464 392638 147520
rect 389270 49544 389326 49600
rect 395710 347112 395766 347168
rect 398378 452104 398434 452160
rect 398102 247152 398158 247208
rect 401506 451424 401562 451480
rect 402518 249600 402574 249656
rect 402426 247968 402482 248024
rect 402610 247696 402666 247752
rect 403806 456048 403862 456104
rect 403990 248104 404046 248160
rect 405094 458904 405150 458960
rect 405186 452920 405242 452976
rect 405002 47912 405058 47968
rect 406198 347384 406254 347440
rect 416778 535880 416834 535936
rect 417054 533704 417110 533760
rect 406842 457544 406898 457600
rect 406658 457408 406714 457464
rect 406474 457136 406530 457192
rect 406382 454008 406438 454064
rect 405462 249736 405518 249792
rect 405278 247832 405334 247888
rect 406750 455640 406806 455696
rect 406934 452784 406990 452840
rect 406842 149232 406898 149288
rect 405186 47776 405242 47832
rect 407762 49408 407818 49464
rect 410522 462440 410578 462496
rect 408314 458768 408370 458824
rect 408130 458360 408186 458416
rect 408222 453056 408278 453112
rect 409142 457272 409198 457328
rect 408130 49272 408186 49328
rect 413282 462576 413338 462632
rect 410706 49544 410762 49600
rect 410890 455912 410946 455968
rect 410982 453192 411038 453248
rect 410982 349152 411038 349208
rect 411902 450064 411958 450120
rect 418066 532788 418068 532808
rect 418068 532788 418120 532808
rect 418120 532788 418122 532808
rect 418066 532752 418122 532788
rect 417698 530984 417754 531040
rect 417422 529896 417478 529952
rect 417698 528128 417754 528184
rect 417606 509904 417662 509960
rect 418066 508272 418122 508328
rect 416778 508000 416834 508056
rect 413466 458224 413522 458280
rect 413558 456864 413614 456920
rect 413650 455776 413706 455832
rect 414478 247560 414534 247616
rect 415214 451560 415270 451616
rect 415122 449928 415178 449984
rect 414938 149096 414994 149152
rect 415858 451968 415914 452024
rect 415858 346296 415914 346352
rect 416594 451832 416650 451888
rect 416410 451696 416466 451752
rect 416226 47232 416282 47288
rect 416410 47096 416466 47152
rect 416778 382744 416834 382800
rect 416870 380976 416926 381032
rect 416778 379888 416834 379944
rect 416778 378120 416834 378176
rect 417330 386824 417386 386880
rect 417238 386280 417294 386336
rect 417238 385872 417294 385928
rect 417146 358264 417202 358320
rect 416962 357992 417018 358048
rect 417054 285640 417110 285696
rect 416870 281016 416926 281072
rect 417698 386824 417754 386880
rect 417606 386280 417662 386336
rect 417882 383696 417938 383752
rect 417514 382744 417570 382800
rect 417790 380976 417846 381032
rect 417698 379888 417754 379944
rect 417606 378120 417662 378176
rect 417330 286864 417386 286920
rect 417238 285912 417294 285968
rect 417238 285640 417294 285696
rect 417238 283736 417294 283792
rect 417054 185952 417110 186008
rect 416870 182008 416926 182064
rect 417422 282784 417478 282840
rect 417330 186904 417386 186960
rect 417238 183776 417294 183832
rect 551006 585148 551008 585168
rect 551008 585148 551060 585168
rect 551060 585148 551062 585168
rect 551006 585112 551062 585148
rect 441618 498072 441674 498128
rect 444378 498072 444434 498128
rect 448518 498072 448574 498128
rect 451278 498072 451334 498128
rect 454682 498072 454738 498128
rect 473358 498072 473414 498128
rect 436190 497256 436246 497312
rect 436098 497120 436154 497176
rect 437478 496848 437534 496904
rect 438858 496848 438914 496904
rect 440238 496848 440294 496904
rect 418066 358264 418122 358320
rect 417882 283736 417938 283792
rect 417790 281016 417846 281072
rect 417698 279928 417754 279984
rect 417606 278704 417662 278760
rect 417422 182824 417478 182880
rect 417238 182008 417294 182064
rect 417238 181056 417294 181112
rect 417054 85856 417110 85912
rect 417238 80960 417294 81016
rect 416778 57976 416834 58032
rect 417882 258032 417938 258088
rect 417790 247560 417846 247616
rect 417514 179968 417570 180024
rect 417514 179424 417570 179480
rect 417606 158344 417662 158400
rect 417422 82864 417478 82920
rect 417698 158108 417700 158128
rect 417700 158108 417752 158128
rect 417752 158108 417754 158128
rect 417698 158072 417754 158108
rect 417606 58248 417662 58304
rect 418618 346296 418674 346352
rect 418618 345616 418674 345672
rect 418618 258304 418674 258360
rect 418342 249464 418398 249520
rect 417882 186904 417938 186960
rect 417790 146920 417846 146976
rect 417974 183776 418030 183832
rect 417882 86808 417938 86864
rect 442998 496984 443054 497040
rect 443090 496848 443146 496904
rect 447138 496984 447194 497040
rect 445758 496848 445814 496904
rect 447230 496848 447286 496904
rect 449990 496984 450046 497040
rect 449898 496848 449954 496904
rect 452658 497528 452714 497584
rect 451370 496848 451426 496904
rect 452750 496848 452806 496904
rect 454038 496848 454094 496904
rect 455418 497120 455474 497176
rect 480350 498092 480406 498128
rect 480350 498072 480352 498092
rect 480352 498072 480404 498092
rect 480404 498072 480406 498092
rect 456890 496984 456946 497040
rect 456798 496848 456854 496904
rect 458270 496984 458326 497040
rect 459558 497004 459614 497040
rect 459558 496984 459560 497004
rect 459560 496984 459612 497004
rect 459612 496984 459614 497004
rect 458178 496848 458234 496904
rect 470782 496984 470838 497040
rect 476118 497004 476174 497040
rect 476118 496984 476120 497004
rect 476120 496984 476172 497004
rect 476172 496984 476174 497004
rect 460938 496848 460994 496904
rect 462318 496848 462374 496904
rect 465078 496848 465134 496904
rect 467838 496848 467894 496904
rect 485778 497936 485834 497992
rect 483018 497120 483074 497176
rect 477498 496868 477554 496904
rect 477498 496848 477500 496868
rect 477500 496848 477552 496868
rect 477552 496848 477554 496868
rect 419630 452648 419686 452704
rect 418066 147056 418122 147112
rect 418986 235864 419042 235920
rect 418618 235456 418674 235512
rect 419170 235592 419226 235648
rect 418710 147056 418766 147112
rect 417974 83680 418030 83736
rect 418802 146920 418858 146976
rect 419538 347828 419540 347848
rect 419540 347828 419592 347848
rect 419592 347828 419594 347848
rect 419538 347792 419594 347828
rect 419998 449792 420054 449848
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 558918 578584 558974 578640
rect 558182 456184 558238 456240
rect 557538 433472 557594 433528
rect 478510 349832 478566 349888
rect 483478 349832 483534 349888
rect 485962 349832 486018 349888
rect 492586 349852 492642 349888
rect 492586 349832 492588 349852
rect 492588 349832 492640 349852
rect 492640 349832 492642 349852
rect 452566 349696 452622 349752
rect 436098 347656 436154 347712
rect 437018 347656 437074 347712
rect 438030 347656 438086 347712
rect 439594 347656 439650 347712
rect 440514 347656 440570 347712
rect 441618 347656 441674 347712
rect 443090 347656 443146 347712
rect 444194 347656 444250 347712
rect 445298 347656 445354 347712
rect 446402 347656 446458 347712
rect 447138 347656 447194 347712
rect 448242 347656 448298 347712
rect 448518 347656 448574 347712
rect 449898 347656 449954 347712
rect 450634 347656 450690 347712
rect 451370 347656 451426 347712
rect 419630 347248 419686 347304
rect 419814 346876 419816 346896
rect 419816 346876 419868 346896
rect 419868 346876 419870 346896
rect 419814 346840 419870 346876
rect 438858 345616 438914 345672
rect 488262 349696 488318 349752
rect 491022 349696 491078 349752
rect 508502 349696 508558 349752
rect 520922 349696 520978 349752
rect 505926 349560 505982 349616
rect 498474 349016 498530 349072
rect 500958 349016 501014 349072
rect 503442 349016 503498 349072
rect 515862 349560 515918 349616
rect 510986 349016 511042 349072
rect 523314 349016 523370 349072
rect 453026 347656 453082 347712
rect 453578 347656 453634 347712
rect 455234 347656 455290 347712
rect 455786 347656 455842 347712
rect 456154 347656 456210 347712
rect 456982 347656 457038 347712
rect 458086 347656 458142 347712
rect 458362 347676 458418 347712
rect 458362 347656 458364 347676
rect 458364 347656 458416 347676
rect 458416 347656 458418 347676
rect 459466 347692 459468 347712
rect 459468 347692 459520 347712
rect 459520 347692 459522 347712
rect 459466 347656 459522 347692
rect 460938 347656 460994 347712
rect 461490 347656 461546 347712
rect 460570 346976 460626 347032
rect 462778 347656 462834 347712
rect 463514 347656 463570 347712
rect 463882 347656 463938 347712
rect 465170 347656 465226 347712
rect 465722 347656 465778 347712
rect 467378 347656 467434 347712
rect 468666 347656 468722 347712
rect 469770 347656 469826 347712
rect 471242 347656 471298 347712
rect 472070 347656 472126 347712
rect 473358 347656 473414 347712
rect 474370 347656 474426 347712
rect 475658 347676 475714 347712
rect 475658 347656 475660 347676
rect 475660 347656 475712 347676
rect 475712 347656 475714 347676
rect 465262 346976 465318 347032
rect 467930 347520 467986 347576
rect 476946 347656 477002 347712
rect 478050 347692 478052 347712
rect 478052 347692 478104 347712
rect 478104 347692 478106 347712
rect 478050 347656 478106 347692
rect 479154 347676 479210 347712
rect 479154 347656 479156 347676
rect 479156 347656 479208 347676
rect 479208 347656 479210 347676
rect 513378 347656 513434 347712
rect 518346 347656 518402 347712
rect 525890 347656 525946 347712
rect 580262 577632 580318 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 558918 429664 558974 429720
rect 551006 335452 551008 335472
rect 551008 335452 551060 335472
rect 551060 335452 551062 335472
rect 551006 335416 551062 335452
rect 485962 249756 486018 249792
rect 485962 249736 485964 249756
rect 485964 249736 486016 249756
rect 486016 249736 486018 249756
rect 488262 249736 488318 249792
rect 491022 249736 491078 249792
rect 495898 249736 495954 249792
rect 498474 249736 498530 249792
rect 500958 249736 501014 249792
rect 503534 249736 503590 249792
rect 470966 249600 471022 249656
rect 483478 249600 483534 249656
rect 473634 249328 473690 249384
rect 505926 249600 505982 249656
rect 508502 249600 508558 249656
rect 515862 249600 515918 249656
rect 520922 249600 520978 249656
rect 443182 248240 443238 248296
rect 447138 248240 447194 248296
rect 449806 248240 449862 248296
rect 436098 247288 436154 247344
rect 436190 247016 436246 247072
rect 437478 247016 437534 247072
rect 438858 247016 438914 247072
rect 440238 247016 440294 247072
rect 441618 247016 441674 247072
rect 444286 247016 444342 247072
rect 441618 235864 441674 235920
rect 440238 235728 440294 235784
rect 438858 235592 438914 235648
rect 437478 235456 437534 235512
rect 445666 247016 445722 247072
rect 447046 247016 447102 247072
rect 450174 248240 450230 248296
rect 450358 248240 450414 248296
rect 451370 248240 451426 248296
rect 452658 248260 452714 248296
rect 452658 248240 452660 248260
rect 452660 248240 452712 248260
rect 452712 248240 452714 248260
rect 448426 247016 448482 247072
rect 455418 248276 455420 248296
rect 455420 248276 455472 248296
rect 455472 248276 455474 248296
rect 455418 248240 455474 248276
rect 462318 248240 462374 248296
rect 467838 248240 467894 248296
rect 460938 247968 460994 248024
rect 461122 247988 461178 248024
rect 461122 247968 461124 247988
rect 461124 247968 461176 247988
rect 461176 247968 461178 247988
rect 465078 247968 465134 248024
rect 461122 247832 461178 247888
rect 463698 247832 463754 247888
rect 469218 247852 469274 247888
rect 469218 247832 469220 247852
rect 469220 247832 469272 247852
rect 469272 247832 469274 247852
rect 455878 247560 455934 247616
rect 462226 247560 462282 247616
rect 452566 247016 452622 247072
rect 457994 247424 458050 247480
rect 453946 247016 454002 247072
rect 455326 247016 455382 247072
rect 458086 247016 458142 247072
rect 473358 247832 473414 247888
rect 466458 247696 466514 247752
rect 478878 247716 478934 247752
rect 478878 247696 478880 247716
rect 478880 247696 478932 247716
rect 478932 247696 478934 247716
rect 465078 247580 465134 247616
rect 465078 247560 465080 247580
rect 465080 247560 465132 247580
rect 465132 247560 465134 247580
rect 470782 247560 470838 247616
rect 476118 247444 476174 247480
rect 476118 247424 476120 247444
rect 476120 247424 476172 247444
rect 476172 247424 476174 247444
rect 459466 247288 459522 247344
rect 471978 247288 472034 247344
rect 473358 247288 473414 247344
rect 477498 247308 477554 247344
rect 477498 247288 477500 247308
rect 477500 247288 477552 247308
rect 477552 247288 477554 247308
rect 480534 247016 480590 247072
rect 492678 247016 492734 247072
rect 510618 247016 510674 247072
rect 513378 247016 513434 247072
rect 523038 247016 523094 247072
rect 525798 247036 525854 247072
rect 525798 247016 525800 247036
rect 525800 247016 525852 247036
rect 525852 247016 525854 247036
rect 459558 238584 459614 238640
rect 558918 329160 558974 329216
rect 550822 235048 550878 235104
rect 458086 149776 458142 149832
rect 478510 149776 478566 149832
rect 480902 149776 480958 149832
rect 483478 149776 483534 149832
rect 485962 149776 486018 149832
rect 440054 149640 440110 149696
rect 438214 149504 438270 149560
rect 436098 147600 436154 147656
rect 437018 147600 437074 147656
rect 437938 147600 437994 147656
rect 430578 146784 430634 146840
rect 439594 147600 439650 147656
rect 456798 149504 456854 149560
rect 443090 147600 443146 147656
rect 444194 147600 444250 147656
rect 445298 147600 445354 147656
rect 446402 147600 446458 147656
rect 447138 147600 447194 147656
rect 448242 147600 448298 147656
rect 448518 147600 448574 147656
rect 449898 147600 449954 147656
rect 450634 147600 450690 147656
rect 451278 147600 451334 147656
rect 452566 147600 452622 147656
rect 453394 147600 453450 147656
rect 453578 147600 453634 147656
rect 454590 147600 454646 147656
rect 455970 147600 456026 147656
rect 440054 147192 440110 147248
rect 440238 147228 440240 147248
rect 440240 147228 440292 147248
rect 440292 147228 440294 147248
rect 440238 147192 440294 147228
rect 463514 149504 463570 149560
rect 465998 149504 466054 149560
rect 468298 149504 468354 149560
rect 470966 149504 471022 149560
rect 459466 148688 459522 148744
rect 459466 148280 459522 148336
rect 458362 147620 458418 147656
rect 488262 149640 488318 149696
rect 491022 149640 491078 149696
rect 495898 149640 495954 149696
rect 503534 149640 503590 149696
rect 505926 149504 505982 149560
rect 508502 149504 508558 149560
rect 510986 149504 511042 149560
rect 515862 149504 515918 149560
rect 518438 149504 518494 149560
rect 513378 148960 513434 149016
rect 520922 148960 520978 149016
rect 523314 148960 523370 149016
rect 525890 148960 525946 149016
rect 458362 147600 458364 147620
rect 458364 147600 458416 147620
rect 458416 147600 458418 147620
rect 461674 147600 461730 147656
rect 462778 147600 462834 147656
rect 463882 147600 463938 147656
rect 465170 147600 465226 147656
rect 466274 147600 466330 147656
rect 467562 147600 467618 147656
rect 468666 147600 468722 147656
rect 469770 147600 469826 147656
rect 471058 147600 471114 147656
rect 472162 147600 472218 147656
rect 473358 147600 473414 147656
rect 474094 147600 474150 147656
rect 476946 147600 477002 147656
rect 478050 147620 478106 147656
rect 478050 147600 478052 147620
rect 478052 147600 478104 147620
rect 478104 147600 478106 147620
rect 557630 229200 557686 229256
rect 551926 136448 551982 136504
rect 456982 49816 457038 49872
rect 458086 49852 458088 49872
rect 458088 49852 458140 49872
rect 458140 49852 458142 49872
rect 458086 49816 458142 49852
rect 478510 49836 478566 49872
rect 478510 49816 478512 49836
rect 478512 49816 478564 49836
rect 478564 49816 478566 49836
rect 436098 48184 436154 48240
rect 437018 48184 437074 48240
rect 438122 48184 438178 48240
rect 439594 48184 439650 48240
rect 443090 48184 443146 48240
rect 444286 48184 444342 48240
rect 448242 48204 448298 48240
rect 448242 48184 448244 48204
rect 448244 48184 448296 48204
rect 448296 48184 448298 48204
rect 450634 48184 450690 48240
rect 453578 48184 453634 48240
rect 454590 48184 454646 48240
rect 455878 48184 455934 48240
rect 445298 48048 445354 48104
rect 446402 48048 446458 48104
rect 449530 48048 449586 48104
rect 447506 47504 447562 47560
rect 452290 48048 452346 48104
rect 453946 48048 454002 48104
rect 450082 47368 450138 47424
rect 450450 47368 450506 47424
rect 451278 47404 451280 47424
rect 451280 47404 451332 47424
rect 451332 47404 451334 47424
rect 451278 47368 451334 47404
rect 480902 49816 480958 49872
rect 473358 49680 473414 49736
rect 488262 49680 488318 49736
rect 495898 49700 495954 49736
rect 495898 49680 495900 49700
rect 495900 49680 495952 49700
rect 495952 49680 495954 49700
rect 459466 49000 459522 49056
rect 458362 48220 458364 48240
rect 458364 48220 458416 48240
rect 458416 48220 458418 48240
rect 458362 48184 458418 48220
rect 456982 48048 457038 48104
rect 461674 48184 461730 48240
rect 462778 48184 462834 48240
rect 463514 48184 463570 48240
rect 463882 48184 463938 48240
rect 465170 48184 465226 48240
rect 465906 48184 465962 48240
rect 466274 48184 466330 48240
rect 467562 48184 467618 48240
rect 468298 48184 468354 48240
rect 468666 48184 468722 48240
rect 469218 48184 469274 48240
rect 470874 48184 470930 48240
rect 471242 48184 471298 48240
rect 472162 48184 472218 48240
rect 459926 47640 459982 47696
rect 469126 48084 469128 48104
rect 469128 48084 469180 48104
rect 469180 48084 469182 48104
rect 469126 48048 469182 48084
rect 503534 49680 503590 49736
rect 493414 49544 493470 49600
rect 498474 49544 498530 49600
rect 500958 49564 501014 49600
rect 500958 49544 500960 49564
rect 500960 49544 501012 49564
rect 501012 49544 501014 49564
rect 505926 49544 505982 49600
rect 508502 49544 508558 49600
rect 510986 49544 511042 49600
rect 513378 49544 513434 49600
rect 515862 49544 515918 49600
rect 520922 49544 520978 49600
rect 525890 49544 525946 49600
rect 474370 48184 474426 48240
rect 475658 48184 475714 48240
rect 476946 48204 477002 48240
rect 476946 48184 476948 48204
rect 476948 48184 477000 48204
rect 477000 48184 477002 48204
rect 478050 48220 478052 48240
rect 478052 48220 478104 48240
rect 478104 48220 478106 48240
rect 478050 48184 478106 48220
rect 563794 459584 563850 459640
rect 558918 229200 558974 229256
rect 558918 129648 558974 129704
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 579986 454416 580042 454472
rect 579618 325216 579674 325272
rect 580170 454280 580226 454336
rect 580078 431568 580134 431624
rect 580078 418240 580134 418296
rect 580078 404912 580134 404968
rect 580078 378392 580134 378448
rect 580078 351872 580134 351928
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 579618 232328 579674 232384
rect 579986 219000 580042 219056
rect 579618 192480 579674 192536
rect 580078 179152 580134 179208
rect 579618 139340 579620 139360
rect 579620 139340 579672 139360
rect 579672 139340 579674 139360
rect 579618 139304 579674 139340
rect 580630 454144 580686 454200
rect 580814 454824 580870 454880
rect 580722 365064 580778 365120
rect 580814 272176 580870 272232
rect 580630 258848 580686 258904
rect 580538 245520 580594 245576
rect 580446 205672 580502 205728
rect 580538 165824 580594 165880
rect 580354 152632 580410 152688
rect 580262 112784 580318 112840
rect 579710 99456 579766 99512
rect 580170 72936 580226 72992
rect 580906 125976 580962 126032
rect 580446 86128 580502 86184
rect 580354 59608 580410 59664
rect 580170 46280 580226 46336
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 46841 682682 46907 682685
rect 244457 682682 244523 682685
rect 46841 682680 244523 682682
rect 46841 682624 46846 682680
rect 46902 682624 244462 682680
rect 244518 682624 244523 682680
rect 46841 682622 244523 682624
rect 46841 682619 46907 682622
rect 244457 682619 244523 682622
rect 197169 682546 197235 682549
rect 390645 682546 390711 682549
rect 197169 682544 390711 682546
rect 197169 682488 197174 682544
rect 197230 682488 390650 682544
rect 390706 682488 390711 682544
rect 197169 682486 390711 682488
rect 197169 682483 197235 682486
rect 390645 682483 390711 682486
rect 53649 682410 53715 682413
rect 247309 682410 247375 682413
rect 53649 682408 247375 682410
rect 53649 682352 53654 682408
rect 53710 682352 247314 682408
rect 247370 682352 247375 682408
rect 53649 682350 247375 682352
rect 53649 682347 53715 682350
rect 247309 682347 247375 682350
rect 51625 682274 51691 682277
rect 247125 682274 247191 682277
rect 51625 682272 247191 682274
rect 51625 682216 51630 682272
rect 51686 682216 247130 682272
rect 247186 682216 247191 682272
rect 51625 682214 247191 682216
rect 51625 682211 51691 682214
rect 247125 682211 247191 682214
rect 137737 682138 137803 682141
rect 193806 682138 193812 682140
rect 137737 682136 193812 682138
rect 137737 682080 137742 682136
rect 137798 682080 193812 682136
rect 137737 682078 193812 682080
rect 137737 682075 137803 682078
rect 193806 682076 193812 682078
rect 193876 682076 193882 682140
rect 195145 682138 195211 682141
rect 390737 682138 390803 682141
rect 195145 682136 390803 682138
rect 195145 682080 195150 682136
rect 195206 682080 390742 682136
rect 390798 682080 390803 682136
rect 195145 682078 390803 682080
rect 195145 682075 195211 682078
rect 390737 682075 390803 682078
rect 75545 682002 75611 682005
rect 186262 682002 186268 682004
rect 75545 682000 186268 682002
rect 75545 681944 75550 682000
rect 75606 681944 186268 682000
rect 75545 681942 186268 681944
rect 75545 681939 75611 681942
rect 186262 681940 186268 681942
rect 186332 681940 186338 682004
rect 192753 682002 192819 682005
rect 390553 682002 390619 682005
rect 192753 682000 390619 682002
rect 192753 681944 192758 682000
rect 192814 681944 390558 682000
rect 390614 681944 390619 682000
rect 192753 681942 390619 681944
rect 192753 681939 192819 681942
rect 390553 681939 390619 681942
rect 168833 681866 168899 681869
rect 193990 681866 193996 681868
rect 168833 681864 193996 681866
rect 168833 681808 168838 681864
rect 168894 681808 193996 681864
rect 168833 681806 193996 681808
rect 168833 681803 168899 681806
rect 193990 681804 193996 681806
rect 194060 681804 194066 681868
rect 60733 681050 60799 681053
rect 236085 681050 236151 681053
rect 60733 681048 236151 681050
rect 60733 680992 60738 681048
rect 60794 680992 236090 681048
rect 236146 680992 236151 681048
rect 60733 680990 236151 680992
rect 60733 680987 60799 680990
rect 236085 680987 236151 680990
rect 34881 680506 34947 680509
rect 240225 680506 240291 680509
rect 34881 680504 240291 680506
rect 34881 680448 34886 680504
rect 34942 680448 240230 680504
rect 240286 680448 240291 680504
rect 34881 680446 240291 680448
rect 34881 680443 34947 680446
rect 240225 680443 240291 680446
rect 30097 680370 30163 680373
rect 237465 680370 237531 680373
rect 30097 680368 237531 680370
rect 30097 680312 30102 680368
rect 30158 680312 237470 680368
rect 237526 680312 237531 680368
rect 30097 680310 237531 680312
rect 30097 680307 30163 680310
rect 237465 680307 237531 680310
rect 169753 679826 169819 679829
rect 250069 679826 250135 679829
rect 169753 679824 250135 679826
rect 169753 679768 169758 679824
rect 169814 679768 250074 679824
rect 250130 679768 250135 679824
rect 169753 679766 250135 679768
rect 169753 679763 169819 679766
rect 250069 679763 250135 679766
rect 144269 679690 144335 679693
rect 255497 679690 255563 679693
rect 144269 679688 255563 679690
rect 144269 679632 144274 679688
rect 144330 679632 255502 679688
rect 255558 679632 255563 679688
rect 144269 679630 255563 679632
rect 144269 679627 144335 679630
rect 255497 679627 255563 679630
rect 79041 679554 79107 679557
rect 237557 679554 237623 679557
rect 79041 679552 237623 679554
rect 79041 679496 79046 679552
rect 79102 679496 237562 679552
rect 237618 679496 237623 679552
rect 79041 679494 237623 679496
rect 79041 679491 79107 679494
rect 237557 679491 237623 679494
rect 190039 679282 190105 679285
rect 190039 679280 190470 679282
rect 190039 679224 190044 679280
rect 190100 679224 190470 679280
rect 190039 679222 190470 679224
rect 190039 679219 190105 679222
rect 190410 679010 190470 679222
rect 389173 679010 389239 679013
rect 190410 679008 389239 679010
rect 190410 678952 389178 679008
rect 389234 678952 389239 679008
rect 190410 678950 389239 678952
rect 389173 678947 389239 678950
rect 186262 678132 186268 678196
rect 186332 678194 186338 678196
rect 254117 678194 254183 678197
rect 186332 678192 254183 678194
rect 186332 678136 254122 678192
rect 254178 678136 254183 678192
rect 186332 678134 254183 678136
rect 186332 678132 186338 678134
rect 254117 678131 254183 678134
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 551001 585172 551067 585173
rect 550950 585170 550956 585172
rect 550910 585110 550956 585170
rect 551020 585168 551067 585172
rect 551062 585112 551067 585168
rect 550950 585108 550956 585110
rect 551020 585108 551067 585112
rect 551001 585107 551067 585108
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 556570 578642 556630 579190
rect 558913 578642 558979 578645
rect 556570 578640 558979 578642
rect 556570 578584 558918 578640
rect 558974 578584 558979 578640
rect 556570 578582 558979 578584
rect 558913 578579 558979 578582
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect 416773 536890 416839 536893
rect 419398 536890 420072 536924
rect 416773 536888 420072 536890
rect 416773 536832 416778 536888
rect 416834 536864 420072 536888
rect 416834 536832 419458 536864
rect 416773 536830 419458 536832
rect 416773 536827 416839 536830
rect 416773 535938 416839 535941
rect 419398 535938 420072 535972
rect 416773 535936 420072 535938
rect 416773 535880 416778 535936
rect 416834 535912 420072 535936
rect 416834 535880 419458 535912
rect 416773 535878 419458 535880
rect 416773 535875 416839 535878
rect 417049 533762 417115 533765
rect 419398 533762 420072 533796
rect 417049 533760 420072 533762
rect 417049 533704 417054 533760
rect 417110 533736 420072 533760
rect 417110 533704 419458 533736
rect 417049 533702 419458 533704
rect 417049 533699 417115 533702
rect 418061 532810 418127 532813
rect 419398 532810 420072 532844
rect 418061 532808 420072 532810
rect 418061 532752 418066 532808
rect 418122 532784 420072 532808
rect 418122 532752 419458 532784
rect 418061 532750 419458 532752
rect 418061 532747 418127 532750
rect 417693 531042 417759 531045
rect 419398 531042 420072 531076
rect 417693 531040 420072 531042
rect 417693 530984 417698 531040
rect 417754 531016 420072 531040
rect 417754 530984 419458 531016
rect 417693 530982 419458 530984
rect 417693 530979 417759 530982
rect 417417 529954 417483 529957
rect 419398 529954 420072 529988
rect 417417 529952 420072 529954
rect 417417 529896 417422 529952
rect 417478 529928 420072 529952
rect 417478 529896 419458 529928
rect 417417 529894 419458 529896
rect 417417 529891 417483 529894
rect 417693 528186 417759 528189
rect 419398 528186 420072 528220
rect 417693 528184 420072 528186
rect 417693 528128 417698 528184
rect 417754 528160 420072 528184
rect 417754 528128 419458 528160
rect 417693 528126 419458 528128
rect 417693 528123 417759 528126
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 417601 509962 417667 509965
rect 419398 509962 420072 509996
rect 417601 509960 420072 509962
rect 417601 509904 417606 509960
rect 417662 509936 420072 509960
rect 417662 509904 419458 509936
rect 417601 509902 419458 509904
rect 417601 509899 417667 509902
rect 418061 508330 418127 508333
rect 419398 508330 420072 508364
rect 418061 508328 420072 508330
rect 418061 508272 418066 508328
rect 418122 508304 420072 508328
rect 418122 508272 419458 508304
rect 418061 508270 419458 508272
rect 418061 508267 418127 508270
rect 416773 508058 416839 508061
rect 419398 508058 420072 508092
rect 416773 508056 420072 508058
rect 416773 508000 416778 508056
rect 416834 508032 420072 508056
rect 416834 508000 419458 508032
rect 416773 507998 419458 508000
rect 416773 507995 416839 507998
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 441613 498132 441679 498133
rect 441613 498128 441660 498132
rect 441724 498130 441730 498132
rect 444373 498130 444439 498133
rect 445334 498130 445340 498132
rect 441613 498072 441618 498128
rect 441613 498068 441660 498072
rect 441724 498070 441770 498130
rect 444373 498128 445340 498130
rect 444373 498072 444378 498128
rect 444434 498072 445340 498128
rect 444373 498070 445340 498072
rect 441724 498068 441730 498070
rect 441613 498067 441679 498068
rect 444373 498067 444439 498070
rect 445334 498068 445340 498070
rect 445404 498068 445410 498132
rect 448513 498130 448579 498133
rect 448646 498130 448652 498132
rect 448513 498128 448652 498130
rect 448513 498072 448518 498128
rect 448574 498072 448652 498128
rect 448513 498070 448652 498072
rect 448513 498067 448579 498070
rect 448646 498068 448652 498070
rect 448716 498068 448722 498132
rect 451273 498130 451339 498133
rect 452326 498130 452332 498132
rect 451273 498128 452332 498130
rect 451273 498072 451278 498128
rect 451334 498072 452332 498128
rect 451273 498070 452332 498072
rect 451273 498067 451339 498070
rect 452326 498068 452332 498070
rect 452396 498068 452402 498132
rect 454677 498130 454743 498133
rect 456190 498130 456196 498132
rect 454677 498128 456196 498130
rect 454677 498072 454682 498128
rect 454738 498072 456196 498128
rect 454677 498070 456196 498072
rect 454677 498067 454743 498070
rect 456190 498068 456196 498070
rect 456260 498068 456266 498132
rect 473353 498130 473419 498133
rect 473486 498130 473492 498132
rect 473353 498128 473492 498130
rect 473353 498072 473358 498128
rect 473414 498072 473492 498128
rect 473353 498070 473492 498072
rect 473353 498067 473419 498070
rect 473486 498068 473492 498070
rect 473556 498068 473562 498132
rect 480345 498130 480411 498133
rect 480846 498130 480852 498132
rect 480345 498128 480852 498130
rect 480345 498072 480350 498128
rect 480406 498072 480852 498128
rect 480345 498070 480852 498072
rect 480345 498067 480411 498070
rect 480846 498068 480852 498070
rect 480916 498068 480922 498132
rect 485773 497994 485839 497997
rect 485998 497994 486004 497996
rect 485773 497992 486004 497994
rect 485773 497936 485778 497992
rect 485834 497936 486004 497992
rect 485773 497934 486004 497936
rect 485773 497931 485839 497934
rect 485998 497932 486004 497934
rect 486068 497932 486074 497996
rect 583520 497844 584960 498084
rect 452653 497586 452719 497589
rect 453430 497586 453436 497588
rect 452653 497584 453436 497586
rect 452653 497528 452658 497584
rect 452714 497528 453436 497584
rect 452653 497526 453436 497528
rect 452653 497523 452719 497526
rect 453430 497524 453436 497526
rect 453500 497524 453506 497588
rect 436185 497314 436251 497317
rect 437054 497314 437060 497316
rect 436185 497312 437060 497314
rect 436185 497256 436190 497312
rect 436246 497256 437060 497312
rect 436185 497254 437060 497256
rect 436185 497251 436251 497254
rect 437054 497252 437060 497254
rect 437124 497252 437130 497316
rect 436093 497180 436159 497181
rect 436093 497178 436140 497180
rect 436048 497176 436140 497178
rect 436048 497120 436098 497176
rect 436048 497118 436140 497120
rect 436093 497116 436140 497118
rect 436204 497116 436210 497180
rect 455413 497178 455479 497181
rect 455822 497178 455828 497180
rect 455413 497176 455828 497178
rect 455413 497120 455418 497176
rect 455474 497120 455828 497176
rect 455413 497118 455828 497120
rect 436093 497115 436159 497116
rect 455413 497115 455479 497118
rect 455822 497116 455828 497118
rect 455892 497116 455898 497180
rect 483013 497178 483079 497181
rect 483422 497178 483428 497180
rect 483013 497176 483428 497178
rect 483013 497120 483018 497176
rect 483074 497120 483428 497176
rect 483013 497118 483428 497120
rect 483013 497115 483079 497118
rect 483422 497116 483428 497118
rect 483492 497116 483498 497180
rect 442993 497042 443059 497045
rect 444230 497042 444236 497044
rect 442993 497040 444236 497042
rect 442993 496984 442998 497040
rect 443054 496984 444236 497040
rect 442993 496982 444236 496984
rect 442993 496979 443059 496982
rect 444230 496980 444236 496982
rect 444300 496980 444306 497044
rect 447133 497042 447199 497045
rect 448278 497042 448284 497044
rect 447133 497040 448284 497042
rect 447133 496984 447138 497040
rect 447194 496984 448284 497040
rect 447133 496982 448284 496984
rect 447133 496979 447199 496982
rect 448278 496980 448284 496982
rect 448348 496980 448354 497044
rect 449985 497042 450051 497045
rect 456885 497044 456951 497045
rect 450670 497042 450676 497044
rect 449985 497040 450676 497042
rect 449985 496984 449990 497040
rect 450046 496984 450676 497040
rect 449985 496982 450676 496984
rect 449985 496979 450051 496982
rect 450670 496980 450676 496982
rect 450740 496980 450746 497044
rect 456885 497042 456932 497044
rect 456840 497040 456932 497042
rect 456840 496984 456890 497040
rect 456840 496982 456932 496984
rect 456885 496980 456932 496982
rect 456996 496980 457002 497044
rect 458265 497042 458331 497045
rect 459318 497042 459324 497044
rect 458265 497040 459324 497042
rect 458265 496984 458270 497040
rect 458326 496984 459324 497040
rect 458265 496982 459324 496984
rect 456885 496979 456951 496980
rect 458265 496979 458331 496982
rect 459318 496980 459324 496982
rect 459388 496980 459394 497044
rect 459553 497042 459619 497045
rect 460606 497042 460612 497044
rect 459553 497040 460612 497042
rect 459553 496984 459558 497040
rect 459614 496984 460612 497040
rect 459553 496982 460612 496984
rect 459553 496979 459619 496982
rect 460606 496980 460612 496982
rect 460676 496980 460682 497044
rect 470777 497042 470843 497045
rect 476113 497044 476179 497045
rect 470910 497042 470916 497044
rect 470777 497040 470916 497042
rect 470777 496984 470782 497040
rect 470838 496984 470916 497040
rect 470777 496982 470916 496984
rect 470777 496979 470843 496982
rect 470910 496980 470916 496982
rect 470980 496980 470986 497044
rect 476062 496980 476068 497044
rect 476132 497042 476179 497044
rect 476132 497040 476224 497042
rect 476174 496984 476224 497040
rect 476132 496982 476224 496984
rect 476132 496980 476179 496982
rect 476113 496979 476179 496980
rect 437473 496906 437539 496909
rect 438342 496906 438348 496908
rect 437473 496904 438348 496906
rect 437473 496848 437478 496904
rect 437534 496848 438348 496904
rect 437473 496846 438348 496848
rect 437473 496843 437539 496846
rect 438342 496844 438348 496846
rect 438412 496844 438418 496908
rect 438853 496906 438919 496909
rect 439630 496906 439636 496908
rect 438853 496904 439636 496906
rect 438853 496848 438858 496904
rect 438914 496848 439636 496904
rect 438853 496846 439636 496848
rect 438853 496843 438919 496846
rect 439630 496844 439636 496846
rect 439700 496844 439706 496908
rect 440233 496906 440299 496909
rect 443085 496908 443151 496909
rect 440550 496906 440556 496908
rect 440233 496904 440556 496906
rect 440233 496848 440238 496904
rect 440294 496848 440556 496904
rect 440233 496846 440556 496848
rect 440233 496843 440299 496846
rect 440550 496844 440556 496846
rect 440620 496844 440626 496908
rect 443085 496906 443132 496908
rect 443040 496904 443132 496906
rect 443040 496848 443090 496904
rect 443040 496846 443132 496848
rect 443085 496844 443132 496846
rect 443196 496844 443202 496908
rect 445753 496906 445819 496909
rect 446438 496906 446444 496908
rect 445753 496904 446444 496906
rect 445753 496848 445758 496904
rect 445814 496848 446444 496904
rect 445753 496846 446444 496848
rect 443085 496843 443151 496844
rect 445753 496843 445819 496846
rect 446438 496844 446444 496846
rect 446508 496844 446514 496908
rect 447225 496906 447291 496909
rect 449893 496908 449959 496909
rect 447542 496906 447548 496908
rect 447225 496904 447548 496906
rect 447225 496848 447230 496904
rect 447286 496848 447548 496904
rect 447225 496846 447548 496848
rect 447225 496843 447291 496846
rect 447542 496844 447548 496846
rect 447612 496844 447618 496908
rect 449893 496906 449940 496908
rect 449848 496904 449940 496906
rect 449848 496848 449898 496904
rect 449848 496846 449940 496848
rect 449893 496844 449940 496846
rect 450004 496844 450010 496908
rect 451038 496844 451044 496908
rect 451108 496906 451114 496908
rect 451365 496906 451431 496909
rect 451108 496904 451431 496906
rect 451108 496848 451370 496904
rect 451426 496848 451431 496904
rect 451108 496846 451431 496848
rect 451108 496844 451114 496846
rect 449893 496843 449959 496844
rect 451365 496843 451431 496846
rect 452745 496906 452811 496909
rect 453614 496906 453620 496908
rect 452745 496904 453620 496906
rect 452745 496848 452750 496904
rect 452806 496848 453620 496904
rect 452745 496846 453620 496848
rect 452745 496843 452811 496846
rect 453614 496844 453620 496846
rect 453684 496844 453690 496908
rect 454033 496906 454099 496909
rect 454534 496906 454540 496908
rect 454033 496904 454540 496906
rect 454033 496848 454038 496904
rect 454094 496848 454540 496904
rect 454033 496846 454540 496848
rect 454033 496843 454099 496846
rect 454534 496844 454540 496846
rect 454604 496844 454610 496908
rect 456793 496906 456859 496909
rect 458030 496906 458036 496908
rect 456793 496904 458036 496906
rect 456793 496848 456798 496904
rect 456854 496848 458036 496904
rect 456793 496846 458036 496848
rect 456793 496843 456859 496846
rect 458030 496844 458036 496846
rect 458100 496844 458106 496908
rect 458173 496906 458239 496909
rect 460933 496908 460999 496909
rect 458398 496906 458404 496908
rect 458173 496904 458404 496906
rect 458173 496848 458178 496904
rect 458234 496848 458404 496904
rect 458173 496846 458404 496848
rect 458173 496843 458239 496846
rect 458398 496844 458404 496846
rect 458468 496844 458474 496908
rect 460933 496904 460980 496908
rect 461044 496906 461050 496908
rect 462313 496906 462379 496909
rect 463550 496906 463556 496908
rect 460933 496848 460938 496904
rect 460933 496844 460980 496848
rect 461044 496846 461090 496906
rect 462313 496904 463556 496906
rect 462313 496848 462318 496904
rect 462374 496848 463556 496904
rect 462313 496846 463556 496848
rect 461044 496844 461050 496846
rect 460933 496843 460999 496844
rect 462313 496843 462379 496846
rect 463550 496844 463556 496846
rect 463620 496844 463626 496908
rect 465073 496906 465139 496909
rect 465942 496906 465948 496908
rect 465073 496904 465948 496906
rect 465073 496848 465078 496904
rect 465134 496848 465948 496904
rect 465073 496846 465948 496848
rect 465073 496843 465139 496846
rect 465942 496844 465948 496846
rect 466012 496844 466018 496908
rect 467833 496906 467899 496909
rect 468334 496906 468340 496908
rect 467833 496904 468340 496906
rect 467833 496848 467838 496904
rect 467894 496848 468340 496904
rect 467833 496846 468340 496848
rect 467833 496843 467899 496846
rect 468334 496844 468340 496846
rect 468404 496844 468410 496908
rect 477493 496906 477559 496909
rect 478454 496906 478460 496908
rect 477493 496904 478460 496906
rect 477493 496848 477498 496904
rect 477554 496848 478460 496904
rect 477493 496846 478460 496848
rect 477493 496843 477559 496846
rect 478454 496844 478460 496846
rect 478524 496844 478530 496908
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 3366 466516 3372 466580
rect 3436 466578 3442 466580
rect 231853 466578 231919 466581
rect 3436 466576 231919 466578
rect 3436 466520 231858 466576
rect 231914 466520 231919 466576
rect 3436 466518 231919 466520
rect 3436 466516 3442 466518
rect 231853 466515 231919 466518
rect 166625 464130 166691 464133
rect 349153 464130 349219 464133
rect 166625 464128 349219 464130
rect 166625 464072 166630 464128
rect 166686 464072 349158 464128
rect 349214 464072 349219 464128
rect 166625 464070 349219 464072
rect 166625 464067 166691 464070
rect 349153 464067 349219 464070
rect 163589 463994 163655 463997
rect 354673 463994 354739 463997
rect 163589 463992 354739 463994
rect 163589 463936 163594 463992
rect 163650 463936 354678 463992
rect 354734 463936 354739 463992
rect 163589 463934 354739 463936
rect 163589 463931 163655 463934
rect 354673 463931 354739 463934
rect 163957 463858 164023 463861
rect 358813 463858 358879 463861
rect 163957 463856 358879 463858
rect 163957 463800 163962 463856
rect 164018 463800 358818 463856
rect 358874 463800 358879 463856
rect 163957 463798 358879 463800
rect 163957 463795 164023 463798
rect 358813 463795 358879 463798
rect 163773 463722 163839 463725
rect 361573 463722 361639 463725
rect 163773 463720 361639 463722
rect 163773 463664 163778 463720
rect 163834 463664 361578 463720
rect 361634 463664 361639 463720
rect 163773 463662 361639 463664
rect 163773 463659 163839 463662
rect 361573 463659 361639 463662
rect 193990 462844 193996 462908
rect 194060 462906 194066 462908
rect 251541 462906 251607 462909
rect 194060 462904 251607 462906
rect 194060 462848 251546 462904
rect 251602 462848 251607 462904
rect 194060 462846 251607 462848
rect 194060 462844 194066 462846
rect 251541 462843 251607 462846
rect 302417 462770 302483 462773
rect 418654 462770 418660 462772
rect 302417 462768 418660 462770
rect -960 462634 480 462724
rect 302417 462712 302422 462768
rect 302478 462712 418660 462768
rect 302417 462710 418660 462712
rect 302417 462707 302483 462710
rect 418654 462708 418660 462710
rect 418724 462708 418730 462772
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 288709 462634 288775 462637
rect 413277 462634 413343 462637
rect 288709 462632 413343 462634
rect 288709 462576 288714 462632
rect 288770 462576 413282 462632
rect 413338 462576 413343 462632
rect 288709 462574 413343 462576
rect 288709 462571 288775 462574
rect 413277 462571 413343 462574
rect 284293 462498 284359 462501
rect 410517 462498 410583 462501
rect 284293 462496 410583 462498
rect 284293 462440 284298 462496
rect 284354 462440 410522 462496
rect 410578 462440 410583 462496
rect 284293 462438 410583 462440
rect 284293 462435 284359 462438
rect 410517 462435 410583 462438
rect 163497 462362 163563 462365
rect 364333 462362 364399 462365
rect 163497 462360 364399 462362
rect 163497 462304 163502 462360
rect 163558 462304 364338 462360
rect 364394 462304 364399 462360
rect 163497 462302 364399 462304
rect 163497 462299 163563 462302
rect 364333 462299 364399 462302
rect 170397 461546 170463 461549
rect 234797 461546 234863 461549
rect 170397 461544 234863 461546
rect 170397 461488 170402 461544
rect 170458 461488 234802 461544
rect 234858 461488 234863 461544
rect 170397 461486 234863 461488
rect 170397 461483 170463 461486
rect 234797 461483 234863 461486
rect 183001 461410 183067 461413
rect 371233 461410 371299 461413
rect 183001 461408 371299 461410
rect 183001 461352 183006 461408
rect 183062 461352 371238 461408
rect 371294 461352 371299 461408
rect 183001 461350 371299 461352
rect 183001 461347 183067 461350
rect 371233 461347 371299 461350
rect 182817 461274 182883 461277
rect 377029 461274 377095 461277
rect 182817 461272 377095 461274
rect 182817 461216 182822 461272
rect 182878 461216 377034 461272
rect 377090 461216 377095 461272
rect 182817 461214 377095 461216
rect 182817 461211 182883 461214
rect 377029 461211 377095 461214
rect 183185 461138 183251 461141
rect 380985 461138 381051 461141
rect 183185 461136 381051 461138
rect 183185 461080 183190 461136
rect 183246 461080 380990 461136
rect 381046 461080 381051 461136
rect 183185 461078 381051 461080
rect 183185 461075 183251 461078
rect 380985 461075 381051 461078
rect 183369 461002 183435 461005
rect 383653 461002 383719 461005
rect 183369 461000 383719 461002
rect 183369 460944 183374 461000
rect 183430 460944 383658 461000
rect 383714 460944 383719 461000
rect 183369 460942 383719 460944
rect 183369 460939 183435 460942
rect 383653 460939 383719 460942
rect 169109 460186 169175 460189
rect 321093 460186 321159 460189
rect 169109 460184 321159 460186
rect 169109 460128 169114 460184
rect 169170 460128 321098 460184
rect 321154 460128 321159 460184
rect 169109 460126 321159 460128
rect 169109 460123 169175 460126
rect 321093 460123 321159 460126
rect 175181 460050 175247 460053
rect 360285 460050 360351 460053
rect 175181 460048 360351 460050
rect 175181 459992 175186 460048
rect 175242 459992 360290 460048
rect 360346 459992 360351 460048
rect 175181 459990 360351 459992
rect 175181 459987 175247 459990
rect 360285 459987 360351 459990
rect 174445 459914 174511 459917
rect 366357 459914 366423 459917
rect 174445 459912 366423 459914
rect 174445 459856 174450 459912
rect 174506 459856 366362 459912
rect 366418 459856 366423 459912
rect 174445 459854 366423 459856
rect 174445 459851 174511 459854
rect 366357 459851 366423 459854
rect 174997 459778 175063 459781
rect 372245 459778 372311 459781
rect 174997 459776 372311 459778
rect 174997 459720 175002 459776
rect 175058 459720 372250 459776
rect 372306 459720 372311 459776
rect 174997 459718 372311 459720
rect 174997 459715 175063 459718
rect 372245 459715 372311 459718
rect 203333 459642 203399 459645
rect 563789 459642 563855 459645
rect 203333 459640 563855 459642
rect 203333 459584 203338 459640
rect 203394 459584 563794 459640
rect 563850 459584 563855 459640
rect 203333 459582 563855 459584
rect 203333 459579 203399 459582
rect 563789 459579 563855 459582
rect 183093 459234 183159 459237
rect 368933 459234 368999 459237
rect 183093 459232 368999 459234
rect 183093 459176 183098 459232
rect 183154 459176 368938 459232
rect 368994 459176 368999 459232
rect 183093 459174 368999 459176
rect 183093 459171 183159 459174
rect 368933 459171 368999 459174
rect 185761 459098 185827 459101
rect 348325 459098 348391 459101
rect 185761 459096 348391 459098
rect 185761 459040 185766 459096
rect 185822 459040 348330 459096
rect 348386 459040 348391 459096
rect 185761 459038 348391 459040
rect 185761 459035 185827 459038
rect 348325 459035 348391 459038
rect 280245 458962 280311 458965
rect 405089 458962 405155 458965
rect 280245 458960 405155 458962
rect 280245 458904 280250 458960
rect 280306 458904 405094 458960
rect 405150 458904 405155 458960
rect 280245 458902 405155 458904
rect 280245 458899 280311 458902
rect 405089 458899 405155 458902
rect 169201 458826 169267 458829
rect 324497 458826 324563 458829
rect 169201 458824 324563 458826
rect 169201 458768 169206 458824
rect 169262 458768 324502 458824
rect 324558 458768 324563 458824
rect 169201 458766 324563 458768
rect 169201 458763 169267 458766
rect 324497 458763 324563 458766
rect 327165 458826 327231 458829
rect 408309 458826 408375 458829
rect 327165 458824 408375 458826
rect 327165 458768 327170 458824
rect 327226 458768 408314 458824
rect 408370 458768 408375 458824
rect 327165 458766 408375 458768
rect 327165 458763 327231 458766
rect 408309 458763 408375 458766
rect 185577 458690 185643 458693
rect 342529 458690 342595 458693
rect 185577 458688 342595 458690
rect 185577 458632 185582 458688
rect 185638 458632 342534 458688
rect 342590 458632 342595 458688
rect 185577 458630 342595 458632
rect 185577 458627 185643 458630
rect 342529 458627 342595 458630
rect 185945 458554 186011 458557
rect 345381 458554 345447 458557
rect 185945 458552 345447 458554
rect 185945 458496 185950 458552
rect 186006 458496 345386 458552
rect 345442 458496 345447 458552
rect 185945 458494 345447 458496
rect 185945 458491 186011 458494
rect 345381 458491 345447 458494
rect 333605 458418 333671 458421
rect 408125 458418 408191 458421
rect 333605 458416 408191 458418
rect 333605 458360 333610 458416
rect 333666 458360 408130 458416
rect 408186 458360 408191 458416
rect 333605 458358 408191 458360
rect 333605 458355 333671 458358
rect 408125 458355 408191 458358
rect 366725 458282 366791 458285
rect 413461 458282 413527 458285
rect 366725 458280 413527 458282
rect 366725 458224 366730 458280
rect 366786 458224 413466 458280
rect 413522 458224 413527 458280
rect 366725 458222 413527 458224
rect 366725 458219 366791 458222
rect 413461 458219 413527 458222
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 180057 457738 180123 457741
rect 309409 457738 309475 457741
rect 180057 457736 309475 457738
rect 180057 457680 180062 457736
rect 180118 457680 309414 457736
rect 309470 457680 309475 457736
rect 180057 457678 309475 457680
rect 180057 457675 180123 457678
rect 309409 457675 309475 457678
rect 300485 457602 300551 457605
rect 406837 457602 406903 457605
rect 300485 457600 406903 457602
rect 300485 457544 300490 457600
rect 300546 457544 406842 457600
rect 406898 457544 406903 457600
rect 300485 457542 406903 457544
rect 300485 457539 300551 457542
rect 406837 457539 406903 457542
rect 193806 457404 193812 457468
rect 193876 457466 193882 457468
rect 255589 457466 255655 457469
rect 193876 457464 255655 457466
rect 193876 457408 255594 457464
rect 255650 457408 255655 457464
rect 193876 457406 255655 457408
rect 193876 457404 193882 457406
rect 255589 457403 255655 457406
rect 292021 457466 292087 457469
rect 406653 457466 406719 457469
rect 292021 457464 406719 457466
rect 292021 457408 292026 457464
rect 292082 457408 406658 457464
rect 406714 457408 406719 457464
rect 292021 457406 406719 457408
rect 292021 457403 292087 457406
rect 406653 457403 406719 457406
rect 287605 457330 287671 457333
rect 409137 457330 409203 457333
rect 287605 457328 409203 457330
rect 287605 457272 287610 457328
rect 287666 457272 409142 457328
rect 409198 457272 409203 457328
rect 287605 457270 409203 457272
rect 287605 457267 287671 457270
rect 409137 457267 409203 457270
rect 182909 457194 182975 457197
rect 289261 457194 289327 457197
rect 182909 457192 289327 457194
rect 182909 457136 182914 457192
rect 182970 457136 289266 457192
rect 289322 457136 289327 457192
rect 182909 457134 289327 457136
rect 182909 457131 182975 457134
rect 289261 457131 289327 457134
rect 296713 457194 296779 457197
rect 406469 457194 406535 457197
rect 296713 457192 406535 457194
rect 296713 457136 296718 457192
rect 296774 457136 406474 457192
rect 406530 457136 406535 457192
rect 296713 457134 406535 457136
rect 296713 457131 296779 457134
rect 406469 457131 406535 457134
rect 188429 457058 188495 457061
rect 326245 457058 326311 457061
rect 188429 457056 326311 457058
rect 188429 457000 188434 457056
rect 188490 457000 326250 457056
rect 326306 457000 326311 457056
rect 188429 456998 326311 457000
rect 188429 456995 188495 456998
rect 326245 456995 326311 456998
rect 188705 456922 188771 456925
rect 332869 456922 332935 456925
rect 188705 456920 332935 456922
rect 188705 456864 188710 456920
rect 188766 456864 332874 456920
rect 332930 456864 332935 456920
rect 188705 456862 332935 456864
rect 188705 456859 188771 456862
rect 332869 456859 332935 456862
rect 357893 456922 357959 456925
rect 413553 456922 413619 456925
rect 357893 456920 413619 456922
rect 357893 456864 357898 456920
rect 357954 456864 413558 456920
rect 413614 456864 413619 456920
rect 357893 456862 413619 456864
rect 357893 456859 357959 456862
rect 413553 456859 413619 456862
rect 157977 456378 158043 456381
rect 365989 456378 366055 456381
rect 157977 456376 366055 456378
rect 157977 456320 157982 456376
rect 158038 456320 365994 456376
rect 366050 456320 366055 456376
rect 157977 456318 366055 456320
rect 157977 456315 158043 456318
rect 365989 456315 366055 456318
rect 202505 456242 202571 456245
rect 558177 456242 558243 456245
rect 202505 456240 558243 456242
rect 202505 456184 202510 456240
rect 202566 456184 558182 456240
rect 558238 456184 558243 456240
rect 202505 456182 558243 456184
rect 202505 456179 202571 456182
rect 558177 456179 558243 456182
rect 163865 456106 163931 456109
rect 285857 456106 285923 456109
rect 163865 456104 285923 456106
rect 163865 456048 163870 456104
rect 163926 456048 285862 456104
rect 285918 456048 285923 456104
rect 163865 456046 285923 456048
rect 163865 456043 163931 456046
rect 285857 456043 285923 456046
rect 315573 456106 315639 456109
rect 403801 456106 403867 456109
rect 315573 456104 403867 456106
rect 315573 456048 315578 456104
rect 315634 456048 403806 456104
rect 403862 456048 403867 456104
rect 315573 456046 403867 456048
rect 315573 456043 315639 456046
rect 403801 456043 403867 456046
rect 360837 455970 360903 455973
rect 410885 455970 410951 455973
rect 360837 455968 410951 455970
rect 360837 455912 360842 455968
rect 360898 455912 410890 455968
rect 410946 455912 410951 455968
rect 360837 455910 410951 455912
rect 360837 455907 360903 455910
rect 410885 455907 410951 455910
rect 363781 455834 363847 455837
rect 413645 455834 413711 455837
rect 363781 455832 413711 455834
rect 363781 455776 363786 455832
rect 363842 455776 413650 455832
rect 413706 455776 413711 455832
rect 363781 455774 413711 455776
rect 363781 455771 363847 455774
rect 413645 455771 413711 455774
rect 19190 455636 19196 455700
rect 19260 455698 19266 455700
rect 283005 455698 283071 455701
rect 19260 455696 283071 455698
rect 19260 455640 283010 455696
rect 283066 455640 283071 455696
rect 19260 455638 283071 455640
rect 19260 455636 19266 455638
rect 283005 455635 283071 455638
rect 304809 455698 304875 455701
rect 406745 455698 406811 455701
rect 304809 455696 406811 455698
rect 304809 455640 304814 455696
rect 304870 455640 406750 455696
rect 406806 455640 406811 455696
rect 304809 455638 406811 455640
rect 304809 455635 304875 455638
rect 406745 455635 406811 455638
rect 158161 455562 158227 455565
rect 363229 455562 363295 455565
rect 158161 455560 363295 455562
rect 158161 455504 158166 455560
rect 158222 455504 363234 455560
rect 363290 455504 363295 455560
rect 158161 455502 363295 455504
rect 158161 455499 158227 455502
rect 363229 455499 363295 455502
rect 379513 455562 379579 455565
rect 389265 455562 389331 455565
rect 379513 455560 389331 455562
rect 379513 455504 379518 455560
rect 379574 455504 389270 455560
rect 389326 455504 389331 455560
rect 379513 455502 389331 455504
rect 379513 455499 379579 455502
rect 389265 455499 389331 455502
rect 200665 454882 200731 454885
rect 580809 454882 580875 454885
rect 200665 454880 580875 454882
rect 200665 454824 200670 454880
rect 200726 454824 580814 454880
rect 580870 454824 580875 454880
rect 200665 454822 580875 454824
rect 200665 454819 200731 454822
rect 580809 454819 580875 454822
rect 168005 454746 168071 454749
rect 233877 454746 233943 454749
rect 168005 454744 233943 454746
rect 168005 454688 168010 454744
rect 168066 454688 233882 454744
rect 233938 454688 233943 454744
rect 168005 454686 233943 454688
rect 168005 454683 168071 454686
rect 233877 454683 233943 454686
rect 283189 454610 283255 454613
rect 418102 454610 418108 454612
rect 283189 454608 418108 454610
rect 283189 454552 283194 454608
rect 283250 454552 418108 454608
rect 283189 454550 418108 454552
rect 283189 454547 283255 454550
rect 418102 454548 418108 454550
rect 418172 454548 418178 454612
rect 202137 454474 202203 454477
rect 579981 454474 580047 454477
rect 202137 454472 580047 454474
rect 202137 454416 202142 454472
rect 202198 454416 579986 454472
rect 580042 454416 580047 454472
rect 202137 454414 580047 454416
rect 202137 454411 202203 454414
rect 579981 454411 580047 454414
rect 201401 454338 201467 454341
rect 580165 454338 580231 454341
rect 201401 454336 580231 454338
rect 201401 454280 201406 454336
rect 201462 454280 580170 454336
rect 580226 454280 580231 454336
rect 201401 454278 580231 454280
rect 201401 454275 201467 454278
rect 580165 454275 580231 454278
rect 201033 454202 201099 454205
rect 580625 454202 580691 454205
rect 201033 454200 580691 454202
rect 201033 454144 201038 454200
rect 201094 454144 580630 454200
rect 580686 454144 580691 454200
rect 201033 454142 580691 454144
rect 201033 454139 201099 454142
rect 580625 454139 580691 454142
rect 185853 454066 185919 454069
rect 283925 454066 283991 454069
rect 185853 454064 283991 454066
rect 185853 454008 185858 454064
rect 185914 454008 283930 454064
rect 283986 454008 283991 454064
rect 185853 454006 283991 454008
rect 185853 454003 185919 454006
rect 283925 454003 283991 454006
rect 383469 454066 383535 454069
rect 406377 454066 406443 454069
rect 383469 454064 406443 454066
rect 383469 454008 383474 454064
rect 383530 454008 406382 454064
rect 406438 454008 406443 454064
rect 383469 454006 406443 454008
rect 383469 454003 383535 454006
rect 406377 454003 406443 454006
rect 291929 453522 291995 453525
rect 393957 453522 394023 453525
rect 291929 453520 394023 453522
rect 291929 453464 291934 453520
rect 291990 453464 393962 453520
rect 394018 453464 394023 453520
rect 291929 453462 394023 453464
rect 291929 453459 291995 453462
rect 393957 453459 394023 453462
rect 19006 453324 19012 453388
rect 19076 453386 19082 453388
rect 300393 453386 300459 453389
rect 19076 453384 300459 453386
rect 19076 453328 300398 453384
rect 300454 453328 300459 453384
rect 19076 453326 300459 453328
rect 19076 453324 19082 453326
rect 300393 453323 300459 453326
rect 304441 453386 304507 453389
rect 392669 453386 392735 453389
rect 304441 453384 392735 453386
rect 304441 453328 304446 453384
rect 304502 453328 392674 453384
rect 392730 453328 392735 453384
rect 304441 453326 392735 453328
rect 304441 453323 304507 453326
rect 392669 453323 392735 453326
rect 189717 453250 189783 453253
rect 305545 453250 305611 453253
rect 189717 453248 305611 453250
rect 189717 453192 189722 453248
rect 189778 453192 305550 453248
rect 305606 453192 305611 453248
rect 189717 453190 305611 453192
rect 189717 453187 189783 453190
rect 305545 453187 305611 453190
rect 330937 453250 331003 453253
rect 410977 453250 411043 453253
rect 330937 453248 411043 453250
rect 330937 453192 330942 453248
rect 330998 453192 410982 453248
rect 411038 453192 411043 453248
rect 330937 453190 411043 453192
rect 330937 453187 331003 453190
rect 410977 453187 411043 453190
rect 192334 453052 192340 453116
rect 192404 453114 192410 453116
rect 318425 453114 318491 453117
rect 192404 453112 318491 453114
rect 192404 453056 318430 453112
rect 318486 453056 318491 453112
rect 192404 453054 318491 453056
rect 192404 453052 192410 453054
rect 318425 453051 318491 453054
rect 327625 453114 327691 453117
rect 408217 453114 408283 453117
rect 327625 453112 408283 453114
rect 327625 453056 327630 453112
rect 327686 453056 408222 453112
rect 408278 453056 408283 453112
rect 327625 453054 408283 453056
rect 327625 453051 327691 453054
rect 408217 453051 408283 453054
rect 169569 452978 169635 452981
rect 313641 452978 313707 452981
rect 169569 452976 313707 452978
rect 169569 452920 169574 452976
rect 169630 452920 313646 452976
rect 313702 452920 313707 452976
rect 169569 452918 313707 452920
rect 169569 452915 169635 452918
rect 313641 452915 313707 452918
rect 382181 452978 382247 452981
rect 405181 452978 405247 452981
rect 382181 452976 405247 452978
rect 382181 452920 382186 452976
rect 382242 452920 405186 452976
rect 405242 452920 405247 452976
rect 382181 452918 405247 452920
rect 382181 452915 382247 452918
rect 405181 452915 405247 452918
rect 3601 452842 3667 452845
rect 229001 452842 229067 452845
rect 3601 452840 229067 452842
rect 3601 452784 3606 452840
rect 3662 452784 229006 452840
rect 229062 452784 229067 452840
rect 3601 452782 229067 452784
rect 3601 452779 3667 452782
rect 229001 452779 229067 452782
rect 380249 452842 380315 452845
rect 406929 452842 406995 452845
rect 380249 452840 406995 452842
rect 380249 452784 380254 452840
rect 380310 452784 406934 452840
rect 406990 452784 406995 452840
rect 380249 452782 406995 452784
rect 380249 452779 380315 452782
rect 406929 452779 406995 452782
rect 191598 452644 191604 452708
rect 191668 452706 191674 452708
rect 195145 452706 195211 452709
rect 191668 452704 195211 452706
rect 191668 452648 195150 452704
rect 195206 452648 195211 452704
rect 191668 452646 195211 452648
rect 191668 452644 191674 452646
rect 195145 452643 195211 452646
rect 324313 452706 324379 452709
rect 419625 452706 419691 452709
rect 324313 452704 419691 452706
rect 324313 452648 324318 452704
rect 324374 452648 419630 452704
rect 419686 452648 419691 452704
rect 324313 452646 419691 452648
rect 324313 452643 324379 452646
rect 419625 452643 419691 452646
rect 190269 452434 190335 452437
rect 194777 452434 194843 452437
rect 190269 452432 194843 452434
rect 190269 452376 190274 452432
rect 190330 452376 194782 452432
rect 194838 452376 194843 452432
rect 190269 452374 194843 452376
rect 190269 452371 190335 452374
rect 194777 452371 194843 452374
rect 157885 452298 157951 452301
rect 315113 452298 315179 452301
rect 157885 452296 315179 452298
rect 157885 452240 157890 452296
rect 157946 452240 315118 452296
rect 315174 452240 315179 452296
rect 157885 452238 315179 452240
rect 157885 452235 157951 452238
rect 315113 452235 315179 452238
rect 187509 452162 187575 452165
rect 195881 452162 195947 452165
rect 187509 452160 195947 452162
rect 187509 452104 187514 452160
rect 187570 452104 195886 452160
rect 195942 452104 195947 452160
rect 187509 452102 195947 452104
rect 187509 452099 187575 452102
rect 195881 452099 195947 452102
rect 383561 452162 383627 452165
rect 398373 452162 398439 452165
rect 383561 452160 398439 452162
rect 383561 452104 383566 452160
rect 383622 452104 398378 452160
rect 398434 452104 398439 452160
rect 383561 452102 398439 452104
rect 383561 452099 383627 452102
rect 398373 452099 398439 452102
rect 15101 452026 15167 452029
rect 230105 452026 230171 452029
rect 15101 452024 230171 452026
rect 15101 451968 15106 452024
rect 15162 451968 230110 452024
rect 230166 451968 230171 452024
rect 15101 451966 230171 451968
rect 15101 451963 15167 451966
rect 230105 451963 230171 451966
rect 295241 452026 295307 452029
rect 415853 452026 415919 452029
rect 295241 452024 415919 452026
rect 295241 451968 295246 452024
rect 295302 451968 415858 452024
rect 415914 451968 415919 452024
rect 295241 451966 415919 451968
rect 295241 451963 295307 451966
rect 415853 451963 415919 451966
rect 193213 451890 193279 451893
rect 227897 451890 227963 451893
rect 193213 451888 227963 451890
rect 193213 451832 193218 451888
rect 193274 451832 227902 451888
rect 227958 451832 227963 451888
rect 193213 451830 227963 451832
rect 193213 451827 193279 451830
rect 227897 451827 227963 451830
rect 352281 451890 352347 451893
rect 383469 451890 383535 451893
rect 352281 451888 383535 451890
rect 352281 451832 352286 451888
rect 352342 451832 383474 451888
rect 383530 451832 383535 451888
rect 352281 451830 383535 451832
rect 352281 451827 352347 451830
rect 383469 451827 383535 451830
rect 384665 451890 384731 451893
rect 416589 451890 416655 451893
rect 384665 451888 416655 451890
rect 384665 451832 384670 451888
rect 384726 451832 416594 451888
rect 416650 451832 416655 451888
rect 384665 451830 416655 451832
rect 384665 451827 384731 451830
rect 416589 451827 416655 451830
rect 180701 451754 180767 451757
rect 280153 451754 280219 451757
rect 180701 451752 280219 451754
rect 180701 451696 180706 451752
rect 180762 451696 280158 451752
rect 280214 451696 280219 451752
rect 180701 451694 280219 451696
rect 180701 451691 180767 451694
rect 280153 451691 280219 451694
rect 375833 451754 375899 451757
rect 416405 451754 416471 451757
rect 375833 451752 416471 451754
rect 375833 451696 375838 451752
rect 375894 451696 416410 451752
rect 416466 451696 416471 451752
rect 375833 451694 416471 451696
rect 375833 451691 375899 451694
rect 416405 451691 416471 451694
rect 158529 451618 158595 451621
rect 303337 451618 303403 451621
rect 158529 451616 303403 451618
rect 158529 451560 158534 451616
rect 158590 451560 303342 451616
rect 303398 451560 303403 451616
rect 158529 451558 303403 451560
rect 158529 451555 158595 451558
rect 303337 451555 303403 451558
rect 308489 451618 308555 451621
rect 415209 451618 415275 451621
rect 308489 451616 415275 451618
rect 308489 451560 308494 451616
rect 308550 451560 415214 451616
rect 415270 451560 415275 451616
rect 308489 451558 415275 451560
rect 308489 451555 308555 451558
rect 415209 451555 415275 451558
rect 190361 451482 190427 451485
rect 193673 451482 193739 451485
rect 190361 451480 193739 451482
rect 190361 451424 190366 451480
rect 190422 451424 193678 451480
rect 193734 451424 193739 451480
rect 190361 451422 193739 451424
rect 190361 451419 190427 451422
rect 193673 451419 193739 451422
rect 360009 451482 360075 451485
rect 401501 451482 401567 451485
rect 360009 451480 401567 451482
rect 360009 451424 360014 451480
rect 360070 451424 401506 451480
rect 401562 451424 401567 451480
rect 360009 451422 401567 451424
rect 360009 451419 360075 451422
rect 401501 451419 401567 451422
rect 191097 450938 191163 450941
rect 357341 450938 357407 450941
rect 191097 450936 357407 450938
rect 191097 450880 191102 450936
rect 191158 450880 357346 450936
rect 357402 450880 357407 450936
rect 191097 450878 357407 450880
rect 191097 450875 191163 450878
rect 357341 450875 357407 450878
rect 344921 450802 344987 450805
rect 388437 450802 388503 450805
rect 344921 450800 388503 450802
rect 344921 450744 344926 450800
rect 344982 450744 388442 450800
rect 388498 450744 388503 450800
rect 344921 450742 388503 450744
rect 344921 450739 344987 450742
rect 388437 450739 388503 450742
rect 190177 450666 190243 450669
rect 197813 450666 197879 450669
rect 190177 450664 197879 450666
rect 190177 450608 190182 450664
rect 190238 450608 197818 450664
rect 197874 450608 197879 450664
rect 190177 450606 197879 450608
rect 190177 450603 190243 450606
rect 197813 450603 197879 450606
rect 350809 450666 350875 450669
rect 388621 450666 388687 450669
rect 350809 450664 388687 450666
rect 350809 450608 350814 450664
rect 350870 450608 388626 450664
rect 388682 450608 388687 450664
rect 350809 450606 388687 450608
rect 350809 450603 350875 450606
rect 388621 450603 388687 450606
rect 156781 450530 156847 450533
rect 210417 450530 210483 450533
rect 156781 450528 210483 450530
rect 156781 450472 156786 450528
rect 156842 450472 210422 450528
rect 210478 450472 210483 450528
rect 156781 450470 210483 450472
rect 156781 450467 156847 450470
rect 210417 450467 210483 450470
rect 322841 450530 322907 450533
rect 418838 450530 418844 450532
rect 322841 450528 418844 450530
rect 322841 450472 322846 450528
rect 322902 450472 418844 450528
rect 322841 450470 418844 450472
rect 322841 450467 322907 450470
rect 418838 450468 418844 450470
rect 418908 450468 418914 450532
rect 193990 450332 193996 450396
rect 194060 450394 194066 450396
rect 194133 450394 194199 450397
rect 194060 450392 194199 450394
rect 194060 450336 194138 450392
rect 194194 450336 194199 450392
rect 194060 450334 194199 450336
rect 194060 450332 194066 450334
rect 194133 450331 194199 450334
rect 353753 450394 353819 450397
rect 392577 450394 392643 450397
rect 353753 450392 392643 450394
rect 353753 450336 353758 450392
rect 353814 450336 392582 450392
rect 392638 450336 392643 450392
rect 353753 450334 392643 450336
rect 353753 450331 353819 450334
rect 392577 450331 392643 450334
rect 183461 450258 183527 450261
rect 351545 450258 351611 450261
rect 183461 450256 351611 450258
rect 183461 450200 183466 450256
rect 183522 450200 351550 450256
rect 351606 450200 351611 450256
rect 183461 450198 351611 450200
rect 183461 450195 183527 450198
rect 351545 450195 351611 450198
rect 358721 450258 358787 450261
rect 415894 450258 415900 450260
rect 358721 450256 415900 450258
rect 358721 450200 358726 450256
rect 358782 450200 415900 450256
rect 358721 450198 415900 450200
rect 358721 450195 358787 450198
rect 415894 450196 415900 450198
rect 415964 450196 415970 450260
rect 156597 450122 156663 450125
rect 360193 450122 360259 450125
rect 156597 450120 360259 450122
rect 156597 450064 156602 450120
rect 156658 450064 360198 450120
rect 360254 450064 360259 450120
rect 156597 450062 360259 450064
rect 156597 450059 156663 450062
rect 360193 450059 360259 450062
rect 378777 450122 378843 450125
rect 411897 450122 411963 450125
rect 378777 450120 411963 450122
rect 378777 450064 378782 450120
rect 378838 450064 411902 450120
rect 411958 450064 411963 450120
rect 378777 450062 411963 450064
rect 378777 450059 378843 450062
rect 411897 450059 411963 450062
rect 14733 449986 14799 449989
rect 232313 449986 232379 449989
rect 14733 449984 232379 449986
rect 14733 449928 14738 449984
rect 14794 449928 232318 449984
rect 232374 449928 232379 449984
rect 14733 449926 232379 449928
rect 14733 449923 14799 449926
rect 232313 449923 232379 449926
rect 279049 449986 279115 449989
rect 415117 449986 415183 449989
rect 279049 449984 415183 449986
rect 279049 449928 279054 449984
rect 279110 449928 415122 449984
rect 415178 449928 415183 449984
rect 279049 449926 415183 449928
rect 279049 449923 279115 449926
rect 415117 449923 415183 449926
rect 229737 449850 229803 449853
rect 6870 449848 229803 449850
rect 6870 449792 229742 449848
rect 229798 449792 229803 449848
rect 6870 449790 229803 449792
rect -960 449578 480 449668
rect 3509 449578 3575 449581
rect -960 449576 3575 449578
rect -960 449520 3514 449576
rect 3570 449520 3575 449576
rect -960 449518 3575 449520
rect -960 449428 480 449518
rect 3509 449515 3575 449518
rect 3509 449442 3575 449445
rect 6870 449442 6930 449790
rect 229737 449787 229803 449790
rect 355593 449850 355659 449853
rect 419993 449850 420059 449853
rect 355593 449848 420059 449850
rect 355593 449792 355598 449848
rect 355654 449792 419998 449848
rect 420054 449792 420059 449848
rect 355593 449790 420059 449792
rect 355593 449787 355659 449790
rect 419993 449787 420059 449790
rect 134333 449714 134399 449717
rect 386137 449714 386203 449717
rect 134333 449712 386203 449714
rect 134333 449656 134338 449712
rect 134394 449656 386142 449712
rect 386198 449656 386203 449712
rect 134333 449654 386203 449656
rect 134333 449651 134399 449654
rect 386137 449651 386203 449654
rect 386413 449714 386479 449717
rect 389214 449714 389220 449716
rect 386413 449712 389220 449714
rect 386413 449656 386418 449712
rect 386474 449656 389220 449712
rect 386413 449654 389220 449656
rect 386413 449651 386479 449654
rect 389214 449652 389220 449654
rect 389284 449652 389290 449716
rect 187417 449578 187483 449581
rect 193213 449578 193279 449581
rect 193949 449578 194015 449581
rect 187417 449576 193279 449578
rect 187417 449520 187422 449576
rect 187478 449520 193218 449576
rect 193274 449520 193279 449576
rect 187417 449518 193279 449520
rect 187417 449515 187483 449518
rect 193213 449515 193279 449518
rect 193676 449576 194015 449578
rect 193676 449520 193954 449576
rect 194010 449520 194015 449576
rect 193676 449518 194015 449520
rect 3509 449440 6930 449442
rect 3509 449384 3514 449440
rect 3570 449384 6930 449440
rect 3509 449382 6930 449384
rect 3509 449379 3575 449382
rect 177757 448762 177823 448765
rect 193676 448762 193736 449518
rect 193949 449515 194015 449518
rect 387609 449578 387675 449581
rect 390001 449578 390067 449581
rect 387609 449576 390067 449578
rect 387609 449520 387614 449576
rect 387670 449520 390006 449576
rect 390062 449520 390067 449576
rect 387609 449518 390067 449520
rect 387609 449515 387675 449518
rect 390001 449515 390067 449518
rect 193806 449244 193812 449308
rect 193876 449306 193882 449308
rect 194041 449306 194107 449309
rect 193876 449304 194107 449306
rect 193876 449248 194046 449304
rect 194102 449248 194107 449304
rect 193876 449246 194107 449248
rect 193876 449244 193882 449246
rect 194041 449243 194107 449246
rect 177757 448760 193736 448762
rect 177757 448704 177762 448760
rect 177818 448704 193736 448760
rect 177757 448702 193736 448704
rect 177757 448699 177823 448702
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 150934 435236 150940 435300
rect 151004 435298 151010 435300
rect 151077 435298 151143 435301
rect 151004 435296 151143 435298
rect 151004 435240 151082 435296
rect 151138 435240 151143 435296
rect 151004 435238 151143 435240
rect 151004 435236 151010 435238
rect 151077 435235 151143 435238
rect 550832 433468 550838 433532
rect 550902 433530 550908 433532
rect 557533 433530 557599 433533
rect 550902 433528 557599 433530
rect 550902 433472 557538 433528
rect 557594 433472 557599 433528
rect 550902 433470 557599 433472
rect 550902 433468 550908 433470
rect 557533 433467 557599 433470
rect 580073 431626 580139 431629
rect 583520 431626 584960 431716
rect 580073 431624 584960 431626
rect 580073 431568 580078 431624
rect 580134 431568 584960 431624
rect 580073 431566 584960 431568
rect 580073 431563 580139 431566
rect 583520 431476 584960 431566
rect 558913 429722 558979 429725
rect 556570 429720 558979 429722
rect 556570 429664 558918 429720
rect 558974 429664 558979 429720
rect 556570 429662 558979 429664
rect 158805 429314 158871 429317
rect 157198 429312 158871 429314
rect 157198 429256 158810 429312
rect 158866 429256 158871 429312
rect 157198 429254 158871 429256
rect 157198 429220 157258 429254
rect 158805 429251 158871 429254
rect 156588 429160 157258 429220
rect 556570 429190 556630 429662
rect 558913 429659 558979 429662
rect -960 423602 480 423692
rect 3233 423602 3299 423605
rect -960 423600 3299 423602
rect -960 423544 3238 423600
rect 3294 423544 3299 423600
rect -960 423542 3299 423544
rect -960 423452 480 423542
rect 3233 423539 3299 423542
rect 580073 418298 580139 418301
rect 583520 418298 584960 418388
rect 580073 418296 584960 418298
rect 580073 418240 580078 418296
rect 580134 418240 584960 418296
rect 580073 418238 584960 418240
rect 580073 418235 580139 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580073 404970 580139 404973
rect 583520 404970 584960 405060
rect 580073 404968 584960 404970
rect 580073 404912 580078 404968
rect 580134 404912 584960 404968
rect 580073 404910 584960 404912
rect 580073 404907 580139 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 4061 397490 4127 397493
rect -960 397488 4127 397490
rect -960 397432 4066 397488
rect 4122 397432 4127 397488
rect -960 397430 4127 397432
rect -960 397340 480 397430
rect 4061 397427 4127 397430
rect 583520 391628 584960 391868
rect 19382 386885 20056 386924
rect 17585 386882 17651 386885
rect 19333 386882 20056 386885
rect 17585 386880 20056 386882
rect 17585 386824 17590 386880
rect 17646 386824 19338 386880
rect 19394 386864 20056 386880
rect 417325 386882 417391 386885
rect 417693 386882 417759 386885
rect 419398 386882 420072 386924
rect 417325 386880 420072 386882
rect 19394 386824 19442 386864
rect 17585 386822 19442 386824
rect 417325 386824 417330 386880
rect 417386 386824 417698 386880
rect 417754 386864 420072 386880
rect 417754 386824 419458 386864
rect 417325 386822 419458 386824
rect 17585 386819 17651 386822
rect 19333 386819 19399 386822
rect 417325 386819 417391 386822
rect 417693 386819 417759 386822
rect 417233 386338 417299 386341
rect 417601 386338 417667 386341
rect 417233 386336 417667 386338
rect 417233 386280 417238 386336
rect 417294 386280 417606 386336
rect 417662 386280 417667 386336
rect 417233 386278 417667 386280
rect 417233 386275 417299 386278
rect 417601 386275 417667 386278
rect 17217 385930 17283 385933
rect 18781 385930 18847 385933
rect 19382 385930 20056 385972
rect 17217 385928 20056 385930
rect 17217 385872 17222 385928
rect 17278 385872 18786 385928
rect 18842 385912 20056 385928
rect 417233 385930 417299 385933
rect 419398 385930 420072 385972
rect 417233 385928 420072 385930
rect 18842 385872 19442 385912
rect 17217 385870 19442 385872
rect 417233 385872 417238 385928
rect 417294 385912 420072 385928
rect 417294 385872 419458 385912
rect 417233 385870 419458 385872
rect 17217 385867 17283 385870
rect 18781 385867 18847 385870
rect 417233 385867 417299 385870
rect -960 384284 480 384524
rect 18873 383754 18939 383757
rect 19382 383754 20056 383796
rect 18873 383752 20056 383754
rect 18873 383696 18878 383752
rect 18934 383736 20056 383752
rect 417877 383754 417943 383757
rect 419398 383754 420072 383796
rect 417877 383752 420072 383754
rect 18934 383696 19442 383736
rect 18873 383694 19442 383696
rect 417877 383696 417882 383752
rect 417938 383736 420072 383752
rect 417938 383696 419458 383736
rect 417877 383694 419458 383696
rect 18873 383691 18939 383694
rect 417877 383691 417943 383694
rect 18965 382802 19031 382805
rect 19382 382802 20056 382844
rect 18965 382800 20056 382802
rect 18965 382744 18970 382800
rect 19026 382784 20056 382800
rect 416773 382802 416839 382805
rect 417509 382802 417575 382805
rect 419398 382802 420072 382844
rect 416773 382800 420072 382802
rect 19026 382744 19442 382784
rect 18965 382742 19442 382744
rect 416773 382744 416778 382800
rect 416834 382744 417514 382800
rect 417570 382784 420072 382800
rect 417570 382744 419458 382784
rect 416773 382742 419458 382744
rect 18965 382739 19031 382742
rect 416773 382739 416839 382742
rect 417509 382739 417575 382742
rect 16757 381034 16823 381037
rect 19057 381034 19123 381037
rect 19382 381034 20056 381076
rect 16757 381032 20056 381034
rect 16757 380976 16762 381032
rect 16818 380976 19062 381032
rect 19118 381016 20056 381032
rect 416865 381034 416931 381037
rect 417785 381034 417851 381037
rect 419398 381034 420072 381076
rect 416865 381032 420072 381034
rect 19118 380976 19442 381016
rect 16757 380974 19442 380976
rect 416865 380976 416870 381032
rect 416926 380976 417790 381032
rect 417846 381016 420072 381032
rect 417846 380976 419458 381016
rect 416865 380974 419458 380976
rect 16757 380971 16823 380974
rect 19057 380971 19123 380974
rect 416865 380971 416931 380974
rect 417785 380971 417851 380974
rect 17309 379946 17375 379949
rect 19382 379946 20056 379988
rect 17309 379944 20056 379946
rect 17309 379888 17314 379944
rect 17370 379928 20056 379944
rect 416773 379946 416839 379949
rect 417693 379946 417759 379949
rect 419398 379946 420072 379988
rect 416773 379944 420072 379946
rect 17370 379888 19442 379928
rect 17309 379886 19442 379888
rect 416773 379888 416778 379944
rect 416834 379888 417698 379944
rect 417754 379928 420072 379944
rect 417754 379888 419458 379928
rect 416773 379886 419458 379888
rect 17309 379883 17375 379886
rect 416773 379883 416839 379886
rect 417693 379883 417759 379886
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect 17401 378178 17467 378181
rect 17769 378178 17835 378181
rect 19382 378178 20056 378220
rect 17401 378176 20056 378178
rect 17401 378120 17406 378176
rect 17462 378120 17774 378176
rect 17830 378160 20056 378176
rect 416773 378178 416839 378181
rect 417601 378178 417667 378181
rect 419398 378178 420072 378220
rect 416773 378176 420072 378178
rect 17830 378120 19442 378160
rect 17401 378118 19442 378120
rect 416773 378120 416778 378176
rect 416834 378120 417606 378176
rect 417662 378160 420072 378176
rect 417662 378120 419458 378160
rect 416773 378118 419458 378120
rect 17401 378115 17467 378118
rect 17769 378115 17835 378118
rect 416773 378115 416839 378118
rect 417601 378115 417667 378118
rect -960 371378 480 371468
rect 3969 371378 4035 371381
rect -960 371376 4035 371378
rect -960 371320 3974 371376
rect 4030 371320 4035 371376
rect -960 371318 4035 371320
rect -960 371228 480 371318
rect 3969 371315 4035 371318
rect 580717 365122 580783 365125
rect 583520 365122 584960 365212
rect 580717 365120 584960 365122
rect 580717 365064 580722 365120
rect 580778 365064 584960 365120
rect 580717 365062 584960 365064
rect 580717 365059 580783 365062
rect 583520 364972 584960 365062
rect 16941 359954 17007 359957
rect 19149 359954 19215 359957
rect 19382 359954 20056 359996
rect 417918 359954 417924 359956
rect 16941 359952 20056 359954
rect 16941 359896 16946 359952
rect 17002 359896 19154 359952
rect 19210 359936 20056 359952
rect 19210 359896 19442 359936
rect 16941 359894 19442 359896
rect 412590 359894 417924 359954
rect 16941 359891 17007 359894
rect 19149 359891 19215 359894
rect 390001 359410 390067 359413
rect 412590 359410 412650 359894
rect 417918 359892 417924 359894
rect 417988 359954 417994 359956
rect 419398 359954 420072 359996
rect 417988 359936 420072 359954
rect 417988 359894 419458 359936
rect 417988 359892 417994 359894
rect 390001 359408 412650 359410
rect 390001 359352 390006 359408
rect 390062 359352 412650 359408
rect 390001 359350 412650 359352
rect 390001 359347 390067 359350
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 17033 358322 17099 358325
rect 19382 358322 20056 358364
rect 17033 358320 20056 358322
rect 17033 358264 17038 358320
rect 17094 358304 20056 358320
rect 417141 358322 417207 358325
rect 418061 358322 418127 358325
rect 419398 358322 420072 358364
rect 417141 358320 420072 358322
rect 17094 358264 19442 358304
rect 17033 358262 19442 358264
rect 417141 358264 417146 358320
rect 417202 358264 418066 358320
rect 418122 358304 420072 358320
rect 418122 358264 419458 358304
rect 417141 358262 419458 358264
rect 17033 358259 17099 358262
rect 417141 358259 417207 358262
rect 418061 358259 418127 358262
rect 19241 358050 19307 358053
rect 19750 358050 20056 358092
rect 19241 358048 20056 358050
rect 19241 357992 19246 358048
rect 19302 358032 20056 358048
rect 416957 358050 417023 358053
rect 419398 358050 420072 358092
rect 416957 358048 420072 358050
rect 19302 357992 19810 358032
rect 19241 357990 19810 357992
rect 416957 357992 416962 358048
rect 417018 358032 420072 358048
rect 417018 357992 419458 358032
rect 416957 357990 419458 357992
rect 19241 357987 19307 357990
rect 416957 357987 417023 357990
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect 91001 349892 91067 349893
rect 93485 349892 93551 349893
rect 98545 349892 98611 349893
rect 103513 349892 103579 349893
rect 478505 349892 478571 349893
rect 90992 349890 90998 349892
rect 90910 349830 90998 349890
rect 90992 349828 90998 349830
rect 91062 349828 91068 349892
rect 93440 349890 93446 349892
rect 93394 349830 93446 349890
rect 93510 349888 93551 349892
rect 98472 349890 98478 349892
rect 93546 349832 93551 349888
rect 93440 349828 93446 349830
rect 93510 349828 93551 349832
rect 98454 349830 98478 349890
rect 98472 349828 98478 349830
rect 98542 349888 98611 349892
rect 98542 349832 98550 349888
rect 98606 349832 98611 349888
rect 98542 349828 98611 349832
rect 103504 349828 103510 349892
rect 103574 349890 103580 349892
rect 478480 349890 478486 349892
rect 103574 349830 103666 349890
rect 478414 349830 478486 349890
rect 478550 349888 478571 349892
rect 478566 349832 478571 349888
rect 103574 349828 103580 349830
rect 478480 349828 478486 349830
rect 478550 349828 478571 349832
rect 91001 349827 91067 349828
rect 93485 349827 93551 349828
rect 98545 349827 98611 349828
rect 103513 349827 103579 349828
rect 478505 349827 478571 349828
rect 483473 349892 483539 349893
rect 485957 349892 486023 349893
rect 483473 349888 483518 349892
rect 483582 349890 483588 349892
rect 483473 349832 483478 349888
rect 483473 349828 483518 349832
rect 483582 349830 483630 349890
rect 485957 349888 485966 349892
rect 486030 349890 486036 349892
rect 492581 349890 492647 349893
rect 495888 349890 495894 349892
rect 485957 349832 485962 349888
rect 483582 349828 483588 349830
rect 485957 349828 485966 349832
rect 486030 349830 486114 349890
rect 492581 349888 495894 349890
rect 492581 349832 492586 349888
rect 492642 349832 495894 349888
rect 492581 349830 495894 349832
rect 486030 349828 486036 349830
rect 483473 349827 483539 349828
rect 485957 349827 486023 349828
rect 492581 349827 492647 349830
rect 495888 349828 495894 349830
rect 495958 349828 495964 349892
rect 452368 349692 452374 349756
rect 452438 349754 452444 349756
rect 452561 349754 452627 349757
rect 452438 349752 452627 349754
rect 452438 349696 452566 349752
rect 452622 349696 452627 349752
rect 452438 349694 452627 349696
rect 452438 349692 452444 349694
rect 452561 349691 452627 349694
rect 488257 349756 488323 349757
rect 491017 349756 491083 349757
rect 488257 349752 488278 349756
rect 488342 349754 488348 349756
rect 490992 349754 490998 349756
rect 488257 349696 488262 349752
rect 488257 349692 488278 349696
rect 488342 349694 488414 349754
rect 490926 349694 490998 349754
rect 491062 349752 491083 349756
rect 491078 349696 491083 349752
rect 488342 349692 488348 349694
rect 490992 349692 490998 349694
rect 491062 349692 491083 349696
rect 488257 349691 488323 349692
rect 491017 349691 491083 349692
rect 508497 349756 508563 349757
rect 520917 349756 520983 349757
rect 508497 349752 508542 349756
rect 508606 349754 508612 349756
rect 520912 349754 520918 349756
rect 508497 349696 508502 349752
rect 508497 349692 508542 349696
rect 508606 349694 508654 349754
rect 520826 349694 520918 349754
rect 508606 349692 508612 349694
rect 520912 349692 520918 349694
rect 520982 349692 520988 349756
rect 508497 349691 508563 349692
rect 520917 349691 520983 349692
rect 38224 349556 38230 349620
rect 38294 349618 38300 349620
rect 38469 349618 38535 349621
rect 50797 349620 50863 349621
rect 56041 349620 56107 349621
rect 58525 349620 58591 349621
rect 61101 349620 61167 349621
rect 62849 349620 62915 349621
rect 68737 349620 68803 349621
rect 72233 349620 72299 349621
rect 505921 349620 505987 349621
rect 515857 349620 515923 349621
rect 50736 349618 50742 349620
rect 38294 349616 38535 349618
rect 38294 349560 38474 349616
rect 38530 349560 38535 349616
rect 38294 349558 38535 349560
rect 50706 349558 50742 349618
rect 50806 349616 50863 349620
rect 50858 349560 50863 349616
rect 38294 349556 38300 349558
rect 38469 349555 38535 349558
rect 50736 349556 50742 349558
rect 50806 349556 50863 349560
rect 56040 349556 56046 349620
rect 56110 349618 56116 349620
rect 58488 349618 58494 349620
rect 56110 349558 56198 349618
rect 58434 349558 58494 349618
rect 58558 349616 58591 349620
rect 61072 349618 61078 349620
rect 58586 349560 58591 349616
rect 56110 349556 56116 349558
rect 58488 349556 58494 349558
rect 58558 349556 58591 349560
rect 61010 349558 61078 349618
rect 61142 349616 61167 349620
rect 62840 349618 62846 349620
rect 61162 349560 61167 349616
rect 61072 349556 61078 349558
rect 61142 349556 61167 349560
rect 62758 349558 62846 349618
rect 62840 349556 62846 349558
rect 62910 349556 62916 349620
rect 68688 349618 68694 349620
rect 68646 349558 68694 349618
rect 68758 349616 68803 349620
rect 72224 349618 72230 349620
rect 68798 349560 68803 349616
rect 68688 349556 68694 349558
rect 68758 349556 68803 349560
rect 72142 349558 72230 349618
rect 72224 349556 72230 349558
rect 72294 349556 72300 349620
rect 505921 349616 505958 349620
rect 506022 349618 506028 349620
rect 505921 349560 505926 349616
rect 505921 349556 505958 349560
rect 506022 349558 506078 349618
rect 515857 349616 515886 349620
rect 515950 349618 515956 349620
rect 515857 349560 515862 349616
rect 506022 349556 506028 349558
rect 515857 349556 515886 349560
rect 515950 349558 516014 349618
rect 515950 349556 515956 349558
rect 50797 349555 50863 349556
rect 56041 349555 56107 349556
rect 58525 349555 58591 349556
rect 61101 349555 61167 349556
rect 62849 349555 62915 349556
rect 68737 349555 68803 349556
rect 72233 349555 72299 349556
rect 505921 349555 505987 349556
rect 515857 349555 515923 349556
rect 410977 349210 411043 349213
rect 480846 349210 480852 349212
rect 410977 349208 480852 349210
rect 410977 349152 410982 349208
rect 411038 349152 480852 349208
rect 410977 349150 480852 349152
rect 410977 349147 411043 349150
rect 480846 349148 480852 349150
rect 480916 349148 480922 349212
rect 53649 349076 53715 349077
rect 53598 349074 53604 349076
rect 53558 349014 53604 349074
rect 53668 349072 53715 349076
rect 53710 349016 53715 349072
rect 53598 349012 53604 349014
rect 53668 349012 53715 349016
rect 61878 349012 61884 349076
rect 61948 349074 61954 349076
rect 62021 349074 62087 349077
rect 68369 349076 68435 349077
rect 78489 349076 78555 349077
rect 86033 349076 86099 349077
rect 68318 349074 68324 349076
rect 61948 349072 62087 349074
rect 61948 349016 62026 349072
rect 62082 349016 62087 349072
rect 61948 349014 62087 349016
rect 68278 349014 68324 349074
rect 68388 349072 68435 349076
rect 78438 349074 78444 349076
rect 68430 349016 68435 349072
rect 61948 349012 61954 349014
rect 53649 349011 53715 349012
rect 62021 349011 62087 349014
rect 68318 349012 68324 349014
rect 68388 349012 68435 349016
rect 78398 349014 78444 349074
rect 78508 349072 78555 349076
rect 85982 349074 85988 349076
rect 78550 349016 78555 349072
rect 78438 349012 78444 349014
rect 78508 349012 78555 349016
rect 85942 349014 85988 349074
rect 86052 349072 86099 349076
rect 86094 349016 86099 349072
rect 85982 349012 85988 349014
rect 86052 349012 86099 349016
rect 88190 349012 88196 349076
rect 88260 349074 88266 349076
rect 175089 349074 175155 349077
rect 88260 349072 175155 349074
rect 88260 349016 175094 349072
rect 175150 349016 175155 349072
rect 88260 349014 175155 349016
rect 88260 349012 88266 349014
rect 68369 349011 68435 349012
rect 78489 349011 78555 349012
rect 86033 349011 86099 349012
rect 175089 349011 175155 349014
rect 498469 349076 498535 349077
rect 500953 349076 501019 349077
rect 498469 349072 498516 349076
rect 498580 349074 498586 349076
rect 500902 349074 500908 349076
rect 498469 349016 498474 349072
rect 498469 349012 498516 349016
rect 498580 349014 498626 349074
rect 500862 349014 500908 349074
rect 500972 349072 501019 349076
rect 501014 349016 501019 349072
rect 498580 349012 498586 349014
rect 500902 349012 500908 349014
rect 500972 349012 501019 349016
rect 498469 349011 498535 349012
rect 500953 349011 501019 349012
rect 503437 349076 503503 349077
rect 510981 349076 511047 349077
rect 523309 349076 523375 349077
rect 503437 349072 503484 349076
rect 503548 349074 503554 349076
rect 503437 349016 503442 349072
rect 503437 349012 503484 349016
rect 503548 349014 503594 349074
rect 510981 349072 511028 349076
rect 511092 349074 511098 349076
rect 510981 349016 510986 349072
rect 503548 349012 503554 349014
rect 510981 349012 511028 349016
rect 511092 349014 511138 349074
rect 523309 349072 523356 349076
rect 523420 349074 523426 349076
rect 523309 349016 523314 349072
rect 511092 349012 511098 349014
rect 523309 349012 523356 349016
rect 523420 349014 523466 349074
rect 523420 349012 523426 349014
rect 503437 349011 503503 349012
rect 510981 349011 511047 349012
rect 523309 349011 523375 349012
rect 190821 348666 190887 348669
rect 191741 348666 191807 348669
rect 190821 348664 191807 348666
rect 190821 348608 190826 348664
rect 190882 348608 191746 348664
rect 191802 348608 191807 348664
rect 190821 348606 191807 348608
rect 190821 348603 190887 348606
rect 191741 348603 191807 348606
rect 74349 348532 74415 348533
rect 74349 348528 74396 348532
rect 74460 348530 74466 348532
rect 74349 348472 74354 348528
rect 74349 348468 74396 348472
rect 74460 348470 74506 348530
rect 74460 348468 74466 348470
rect 74349 348467 74415 348468
rect 419533 347850 419599 347853
rect 419758 347850 419764 347852
rect 419533 347848 419764 347850
rect 419533 347792 419538 347848
rect 419594 347792 419764 347848
rect 419533 347790 419764 347792
rect 419533 347787 419599 347790
rect 419758 347788 419764 347790
rect 419828 347788 419834 347852
rect 36169 347716 36235 347717
rect 36118 347714 36124 347716
rect 36078 347654 36124 347714
rect 36188 347712 36235 347716
rect 36230 347656 36235 347712
rect 36118 347652 36124 347654
rect 36188 347652 36235 347656
rect 36169 347651 36235 347652
rect 39573 347716 39639 347717
rect 39573 347712 39620 347716
rect 39684 347714 39690 347716
rect 42793 347714 42859 347717
rect 44173 347716 44239 347717
rect 45369 347716 45435 347717
rect 43110 347714 43116 347716
rect 39573 347656 39578 347712
rect 39573 347652 39620 347656
rect 39684 347654 39730 347714
rect 42793 347712 43116 347714
rect 42793 347656 42798 347712
rect 42854 347656 43116 347712
rect 42793 347654 43116 347656
rect 39684 347652 39690 347654
rect 39573 347651 39639 347652
rect 42793 347651 42859 347654
rect 43110 347652 43116 347654
rect 43180 347652 43186 347716
rect 44173 347712 44220 347716
rect 44284 347714 44290 347716
rect 45318 347714 45324 347716
rect 44173 347656 44178 347712
rect 44173 347652 44220 347656
rect 44284 347654 44330 347714
rect 45278 347654 45324 347714
rect 45388 347712 45435 347716
rect 45430 347656 45435 347712
rect 44284 347652 44290 347654
rect 45318 347652 45324 347654
rect 45388 347652 45435 347656
rect 44173 347651 44239 347652
rect 45369 347651 45435 347652
rect 46565 347716 46631 347717
rect 47577 347716 47643 347717
rect 46565 347712 46612 347716
rect 46676 347714 46682 347716
rect 47526 347714 47532 347716
rect 46565 347656 46570 347712
rect 46565 347652 46612 347656
rect 46676 347654 46722 347714
rect 47486 347654 47532 347714
rect 47596 347712 47643 347716
rect 47638 347656 47643 347712
rect 46676 347652 46682 347654
rect 47526 347652 47532 347654
rect 47596 347652 47643 347656
rect 46565 347651 46631 347652
rect 47577 347651 47643 347652
rect 48589 347716 48655 347717
rect 50061 347716 50127 347717
rect 51257 347716 51323 347717
rect 52361 347716 52427 347717
rect 53465 347716 53531 347717
rect 48589 347712 48636 347716
rect 48700 347714 48706 347716
rect 48589 347656 48594 347712
rect 48589 347652 48636 347656
rect 48700 347654 48746 347714
rect 50061 347712 50108 347716
rect 50172 347714 50178 347716
rect 51206 347714 51212 347716
rect 50061 347656 50066 347712
rect 48700 347652 48706 347654
rect 50061 347652 50108 347656
rect 50172 347654 50218 347714
rect 51166 347654 51212 347714
rect 51276 347712 51323 347716
rect 52310 347714 52316 347716
rect 51318 347656 51323 347712
rect 50172 347652 50178 347654
rect 51206 347652 51212 347654
rect 51276 347652 51323 347656
rect 52270 347654 52316 347714
rect 52380 347712 52427 347716
rect 53414 347714 53420 347716
rect 52422 347656 52427 347712
rect 52310 347652 52316 347654
rect 52380 347652 52427 347656
rect 53374 347654 53420 347714
rect 53484 347712 53531 347716
rect 53526 347656 53531 347712
rect 53414 347652 53420 347654
rect 53484 347652 53531 347656
rect 63534 347652 63540 347716
rect 63604 347714 63610 347716
rect 63677 347714 63743 347717
rect 63604 347712 63743 347714
rect 63604 347656 63682 347712
rect 63738 347656 63743 347712
rect 63604 347654 63743 347656
rect 63604 347652 63610 347654
rect 48589 347651 48655 347652
rect 50061 347651 50127 347652
rect 51257 347651 51323 347652
rect 52361 347651 52427 347652
rect 53465 347651 53531 347652
rect 63677 347651 63743 347654
rect 63902 347652 63908 347716
rect 63972 347714 63978 347716
rect 64781 347714 64847 347717
rect 63972 347712 64847 347714
rect 63972 347656 64786 347712
rect 64842 347656 64847 347712
rect 63972 347654 64847 347656
rect 63972 347652 63978 347654
rect 64781 347651 64847 347654
rect 65149 347716 65215 347717
rect 65977 347716 66043 347717
rect 65149 347712 65196 347716
rect 65260 347714 65266 347716
rect 65926 347714 65932 347716
rect 65149 347656 65154 347712
rect 65149 347652 65196 347656
rect 65260 347654 65306 347714
rect 65886 347654 65932 347714
rect 65996 347712 66043 347716
rect 66038 347656 66043 347712
rect 65260 347652 65266 347654
rect 65926 347652 65932 347654
rect 65996 347652 66043 347656
rect 65149 347651 65215 347652
rect 65977 347651 66043 347652
rect 66253 347716 66319 347717
rect 66253 347712 66300 347716
rect 66364 347714 66370 347716
rect 66253 347656 66258 347712
rect 66253 347652 66300 347656
rect 66364 347654 66410 347714
rect 66364 347652 66370 347654
rect 67582 347652 67588 347716
rect 67652 347714 67658 347716
rect 67725 347714 67791 347717
rect 67652 347712 67791 347714
rect 67652 347656 67730 347712
rect 67786 347656 67791 347712
rect 67652 347654 67791 347656
rect 67652 347652 67658 347654
rect 66253 347651 66319 347652
rect 67725 347651 67791 347654
rect 71129 347714 71195 347717
rect 73245 347716 73311 347717
rect 73705 347716 73771 347717
rect 71262 347714 71268 347716
rect 71129 347712 71268 347714
rect 71129 347656 71134 347712
rect 71190 347656 71268 347712
rect 71129 347654 71268 347656
rect 71129 347651 71195 347654
rect 71262 347652 71268 347654
rect 71332 347652 71338 347716
rect 73245 347712 73292 347716
rect 73356 347714 73362 347716
rect 73654 347714 73660 347716
rect 73245 347656 73250 347712
rect 73245 347652 73292 347656
rect 73356 347654 73402 347714
rect 73614 347654 73660 347714
rect 73724 347712 73771 347716
rect 73766 347656 73771 347712
rect 73356 347652 73362 347654
rect 73654 347652 73660 347654
rect 73724 347652 73771 347656
rect 73245 347651 73311 347652
rect 73705 347651 73771 347652
rect 75453 347714 75519 347717
rect 76097 347716 76163 347717
rect 75678 347714 75684 347716
rect 75453 347712 75684 347714
rect 75453 347656 75458 347712
rect 75514 347656 75684 347712
rect 75453 347654 75684 347656
rect 75453 347651 75519 347654
rect 75678 347652 75684 347654
rect 75748 347652 75754 347716
rect 76046 347714 76052 347716
rect 76006 347654 76052 347714
rect 76116 347712 76163 347716
rect 76158 347656 76163 347712
rect 76046 347652 76052 347654
rect 76116 347652 76163 347656
rect 76097 347651 76163 347652
rect 76741 347714 76807 347717
rect 78029 347716 78095 347717
rect 79133 347716 79199 347717
rect 81065 347716 81131 347717
rect 83641 347716 83707 347717
rect 76966 347714 76972 347716
rect 76741 347712 76972 347714
rect 76741 347656 76746 347712
rect 76802 347656 76972 347712
rect 76741 347654 76972 347656
rect 76741 347651 76807 347654
rect 76966 347652 76972 347654
rect 77036 347652 77042 347716
rect 78029 347712 78076 347716
rect 78140 347714 78146 347716
rect 78029 347656 78034 347712
rect 78029 347652 78076 347656
rect 78140 347654 78186 347714
rect 79133 347712 79180 347716
rect 79244 347714 79250 347716
rect 81014 347714 81020 347716
rect 79133 347656 79138 347712
rect 78140 347652 78146 347654
rect 79133 347652 79180 347656
rect 79244 347654 79290 347714
rect 80974 347654 81020 347714
rect 81084 347712 81131 347716
rect 83590 347714 83596 347716
rect 81126 347656 81131 347712
rect 79244 347652 79250 347654
rect 81014 347652 81020 347654
rect 81084 347652 81131 347656
rect 83550 347654 83596 347714
rect 83660 347712 83707 347716
rect 83702 347656 83707 347712
rect 83590 347652 83596 347654
rect 83660 347652 83707 347656
rect 95918 347652 95924 347716
rect 95988 347714 95994 347716
rect 96061 347714 96127 347717
rect 100937 347716 101003 347717
rect 106089 347716 106155 347717
rect 108665 347716 108731 347717
rect 111057 347716 111123 347717
rect 113449 347716 113515 347717
rect 115841 347716 115907 347717
rect 118601 347716 118667 347717
rect 120993 347716 121059 347717
rect 123385 347716 123451 347717
rect 125961 347716 126027 347717
rect 100886 347714 100892 347716
rect 95988 347712 96127 347714
rect 95988 347656 96066 347712
rect 96122 347656 96127 347712
rect 95988 347654 96127 347656
rect 100846 347654 100892 347714
rect 100956 347712 101003 347716
rect 106038 347714 106044 347716
rect 100998 347656 101003 347712
rect 95988 347652 95994 347654
rect 78029 347651 78095 347652
rect 79133 347651 79199 347652
rect 81065 347651 81131 347652
rect 83641 347651 83707 347652
rect 96061 347651 96127 347654
rect 100886 347652 100892 347654
rect 100956 347652 101003 347656
rect 105998 347654 106044 347714
rect 106108 347712 106155 347716
rect 108614 347714 108620 347716
rect 106150 347656 106155 347712
rect 106038 347652 106044 347654
rect 106108 347652 106155 347656
rect 108574 347654 108620 347714
rect 108684 347712 108731 347716
rect 111006 347714 111012 347716
rect 108726 347656 108731 347712
rect 108614 347652 108620 347654
rect 108684 347652 108731 347656
rect 110966 347654 111012 347714
rect 111076 347712 111123 347716
rect 113398 347714 113404 347716
rect 111118 347656 111123 347712
rect 111006 347652 111012 347654
rect 111076 347652 111123 347656
rect 113358 347654 113404 347714
rect 113468 347712 113515 347716
rect 115790 347714 115796 347716
rect 113510 347656 113515 347712
rect 113398 347652 113404 347654
rect 113468 347652 113515 347656
rect 115750 347654 115796 347714
rect 115860 347712 115907 347716
rect 118550 347714 118556 347716
rect 115902 347656 115907 347712
rect 115790 347652 115796 347654
rect 115860 347652 115907 347656
rect 118510 347654 118556 347714
rect 118620 347712 118667 347716
rect 120942 347714 120948 347716
rect 118662 347656 118667 347712
rect 118550 347652 118556 347654
rect 118620 347652 118667 347656
rect 120902 347654 120948 347714
rect 121012 347712 121059 347716
rect 123334 347714 123340 347716
rect 121054 347656 121059 347712
rect 120942 347652 120948 347654
rect 121012 347652 121059 347656
rect 123294 347654 123340 347714
rect 123404 347712 123451 347716
rect 125910 347714 125916 347716
rect 123446 347656 123451 347712
rect 123334 347652 123340 347654
rect 123404 347652 123451 347656
rect 125870 347654 125916 347714
rect 125980 347712 126027 347716
rect 191649 347714 191715 347717
rect 126022 347656 126027 347712
rect 125910 347652 125916 347654
rect 125980 347652 126027 347656
rect 100937 347651 101003 347652
rect 106089 347651 106155 347652
rect 108665 347651 108731 347652
rect 111057 347651 111123 347652
rect 113449 347651 113515 347652
rect 115841 347651 115907 347652
rect 118601 347651 118667 347652
rect 120993 347651 121059 347652
rect 123385 347651 123451 347652
rect 125961 347651 126027 347652
rect 180750 347712 191715 347714
rect 180750 347656 191654 347712
rect 191710 347656 191715 347712
rect 180750 347654 191715 347656
rect 48262 347516 48268 347580
rect 48332 347578 48338 347580
rect 180750 347578 180810 347654
rect 191649 347651 191715 347654
rect 436093 347716 436159 347717
rect 437013 347716 437079 347717
rect 436093 347712 436140 347716
rect 436204 347714 436210 347716
rect 436093 347656 436098 347712
rect 436093 347652 436140 347656
rect 436204 347654 436250 347714
rect 437013 347712 437060 347716
rect 437124 347714 437130 347716
rect 438025 347714 438091 347717
rect 439589 347716 439655 347717
rect 440509 347716 440575 347717
rect 441613 347716 441679 347717
rect 443085 347716 443151 347717
rect 444189 347716 444255 347717
rect 445293 347716 445359 347717
rect 446397 347716 446463 347717
rect 438158 347714 438164 347716
rect 437013 347656 437018 347712
rect 436204 347652 436210 347654
rect 437013 347652 437060 347656
rect 437124 347654 437170 347714
rect 438025 347712 438164 347714
rect 438025 347656 438030 347712
rect 438086 347656 438164 347712
rect 438025 347654 438164 347656
rect 437124 347652 437130 347654
rect 436093 347651 436159 347652
rect 437013 347651 437079 347652
rect 438025 347651 438091 347654
rect 438158 347652 438164 347654
rect 438228 347652 438234 347716
rect 439589 347712 439636 347716
rect 439700 347714 439706 347716
rect 439589 347656 439594 347712
rect 439589 347652 439636 347656
rect 439700 347654 439746 347714
rect 440509 347712 440556 347716
rect 440620 347714 440626 347716
rect 440509 347656 440514 347712
rect 439700 347652 439706 347654
rect 440509 347652 440556 347656
rect 440620 347654 440666 347714
rect 441613 347712 441660 347716
rect 441724 347714 441730 347716
rect 441613 347656 441618 347712
rect 440620 347652 440626 347654
rect 441613 347652 441660 347656
rect 441724 347654 441770 347714
rect 443085 347712 443132 347716
rect 443196 347714 443202 347716
rect 443085 347656 443090 347712
rect 441724 347652 441730 347654
rect 443085 347652 443132 347656
rect 443196 347654 443242 347714
rect 444189 347712 444236 347716
rect 444300 347714 444306 347716
rect 444189 347656 444194 347712
rect 443196 347652 443202 347654
rect 444189 347652 444236 347656
rect 444300 347654 444346 347714
rect 445293 347712 445340 347716
rect 445404 347714 445410 347716
rect 445293 347656 445298 347712
rect 444300 347652 444306 347654
rect 445293 347652 445340 347656
rect 445404 347654 445450 347714
rect 446397 347712 446444 347716
rect 446508 347714 446514 347716
rect 447133 347714 447199 347717
rect 448237 347716 448303 347717
rect 447542 347714 447548 347716
rect 446397 347656 446402 347712
rect 445404 347652 445410 347654
rect 446397 347652 446444 347656
rect 446508 347654 446554 347714
rect 447133 347712 447548 347714
rect 447133 347656 447138 347712
rect 447194 347656 447548 347712
rect 447133 347654 447548 347656
rect 446508 347652 446514 347654
rect 439589 347651 439655 347652
rect 440509 347651 440575 347652
rect 441613 347651 441679 347652
rect 443085 347651 443151 347652
rect 444189 347651 444255 347652
rect 445293 347651 445359 347652
rect 446397 347651 446463 347652
rect 447133 347651 447199 347654
rect 447542 347652 447548 347654
rect 447612 347652 447618 347716
rect 448237 347712 448284 347716
rect 448348 347714 448354 347716
rect 448513 347714 448579 347717
rect 448646 347714 448652 347716
rect 448237 347656 448242 347712
rect 448237 347652 448284 347656
rect 448348 347654 448394 347714
rect 448513 347712 448652 347714
rect 448513 347656 448518 347712
rect 448574 347656 448652 347712
rect 448513 347654 448652 347656
rect 448348 347652 448354 347654
rect 448237 347651 448303 347652
rect 448513 347651 448579 347654
rect 448646 347652 448652 347654
rect 448716 347652 448722 347716
rect 449893 347714 449959 347717
rect 450629 347716 450695 347717
rect 451365 347716 451431 347717
rect 450118 347714 450124 347716
rect 449893 347712 450124 347714
rect 449893 347656 449898 347712
rect 449954 347656 450124 347712
rect 449893 347654 450124 347656
rect 449893 347651 449959 347654
rect 450118 347652 450124 347654
rect 450188 347652 450194 347716
rect 450629 347712 450676 347716
rect 450740 347714 450746 347716
rect 450629 347656 450634 347712
rect 450629 347652 450676 347656
rect 450740 347654 450786 347714
rect 451365 347712 451412 347716
rect 451476 347714 451482 347716
rect 453021 347714 453087 347717
rect 453573 347716 453639 347717
rect 453430 347714 453436 347716
rect 451365 347656 451370 347712
rect 450740 347652 450746 347654
rect 451365 347652 451412 347656
rect 451476 347654 451522 347714
rect 453021 347712 453436 347714
rect 453021 347656 453026 347712
rect 453082 347656 453436 347712
rect 453021 347654 453436 347656
rect 451476 347652 451482 347654
rect 450629 347651 450695 347652
rect 451365 347651 451431 347652
rect 453021 347651 453087 347654
rect 453430 347652 453436 347654
rect 453500 347652 453506 347716
rect 453573 347712 453620 347716
rect 453684 347714 453690 347716
rect 453573 347656 453578 347712
rect 453573 347652 453620 347656
rect 453684 347654 453730 347714
rect 453684 347652 453690 347654
rect 454534 347652 454540 347716
rect 454604 347714 454610 347716
rect 455229 347714 455295 347717
rect 455781 347716 455847 347717
rect 456149 347716 456215 347717
rect 456977 347716 457043 347717
rect 458081 347716 458147 347717
rect 455781 347714 455828 347716
rect 454604 347712 455295 347714
rect 454604 347656 455234 347712
rect 455290 347656 455295 347712
rect 454604 347654 455295 347656
rect 455736 347712 455828 347714
rect 455736 347656 455786 347712
rect 455736 347654 455828 347656
rect 454604 347652 454610 347654
rect 453573 347651 453639 347652
rect 455229 347651 455295 347654
rect 455781 347652 455828 347654
rect 455892 347652 455898 347716
rect 456149 347712 456196 347716
rect 456260 347714 456266 347716
rect 456926 347714 456932 347716
rect 456149 347656 456154 347712
rect 456149 347652 456196 347656
rect 456260 347654 456306 347714
rect 456886 347654 456932 347714
rect 456996 347712 457043 347716
rect 458030 347714 458036 347716
rect 457038 347656 457043 347712
rect 456260 347652 456266 347654
rect 456926 347652 456932 347654
rect 456996 347652 457043 347656
rect 457990 347654 458036 347714
rect 458100 347712 458147 347716
rect 458142 347656 458147 347712
rect 458030 347652 458036 347654
rect 458100 347652 458147 347656
rect 455781 347651 455847 347652
rect 456149 347651 456215 347652
rect 456977 347651 457043 347652
rect 458081 347651 458147 347652
rect 458357 347716 458423 347717
rect 459461 347716 459527 347717
rect 460933 347716 460999 347717
rect 458357 347712 458404 347716
rect 458468 347714 458474 347716
rect 458357 347656 458362 347712
rect 458357 347652 458404 347656
rect 458468 347654 458514 347714
rect 459461 347712 459508 347716
rect 459572 347714 459578 347716
rect 459461 347656 459466 347712
rect 458468 347652 458474 347654
rect 459461 347652 459508 347656
rect 459572 347654 459618 347714
rect 460933 347712 460980 347716
rect 461044 347714 461050 347716
rect 461485 347714 461551 347717
rect 462773 347716 462839 347717
rect 463509 347716 463575 347717
rect 463877 347716 463943 347717
rect 465165 347716 465231 347717
rect 461710 347714 461716 347716
rect 460933 347656 460938 347712
rect 459572 347652 459578 347654
rect 460933 347652 460980 347656
rect 461044 347654 461090 347714
rect 461485 347712 461716 347714
rect 461485 347656 461490 347712
rect 461546 347656 461716 347712
rect 461485 347654 461716 347656
rect 461044 347652 461050 347654
rect 458357 347651 458423 347652
rect 459461 347651 459527 347652
rect 460933 347651 460999 347652
rect 461485 347651 461551 347654
rect 461710 347652 461716 347654
rect 461780 347652 461786 347716
rect 462773 347712 462820 347716
rect 462884 347714 462890 347716
rect 462773 347656 462778 347712
rect 462773 347652 462820 347656
rect 462884 347654 462930 347714
rect 463509 347712 463556 347716
rect 463620 347714 463626 347716
rect 463509 347656 463514 347712
rect 462884 347652 462890 347654
rect 463509 347652 463556 347656
rect 463620 347654 463666 347714
rect 463877 347712 463924 347716
rect 463988 347714 463994 347716
rect 463877 347656 463882 347712
rect 463620 347652 463626 347654
rect 463877 347652 463924 347656
rect 463988 347654 464034 347714
rect 465165 347712 465212 347716
rect 465276 347714 465282 347716
rect 465717 347714 465783 347717
rect 466310 347714 466316 347716
rect 465165 347656 465170 347712
rect 463988 347652 463994 347654
rect 465165 347652 465212 347656
rect 465276 347654 465322 347714
rect 465717 347712 466316 347714
rect 465717 347656 465722 347712
rect 465778 347656 466316 347712
rect 465717 347654 466316 347656
rect 465276 347652 465282 347654
rect 462773 347651 462839 347652
rect 463509 347651 463575 347652
rect 463877 347651 463943 347652
rect 465165 347651 465231 347652
rect 465717 347651 465783 347654
rect 466310 347652 466316 347654
rect 466380 347652 466386 347716
rect 467373 347714 467439 347717
rect 468661 347716 468727 347717
rect 469765 347716 469831 347717
rect 471237 347716 471303 347717
rect 467598 347714 467604 347716
rect 467373 347712 467604 347714
rect 467373 347656 467378 347712
rect 467434 347656 467604 347712
rect 467373 347654 467604 347656
rect 467373 347651 467439 347654
rect 467598 347652 467604 347654
rect 467668 347652 467674 347716
rect 467790 347654 468586 347714
rect 48332 347518 180810 347578
rect 190821 347578 190887 347581
rect 191281 347578 191347 347581
rect 190821 347576 191347 347578
rect 190821 347520 190826 347576
rect 190882 347520 191286 347576
rect 191342 347520 191347 347576
rect 190821 347518 191347 347520
rect 48332 347516 48338 347518
rect 190821 347515 190887 347518
rect 191281 347515 191347 347518
rect 388529 347578 388595 347581
rect 467790 347578 467850 347654
rect 388529 347576 467850 347578
rect 388529 347520 388534 347576
rect 388590 347520 467850 347576
rect 388529 347518 467850 347520
rect 467925 347578 467991 347581
rect 468334 347578 468340 347580
rect 467925 347576 468340 347578
rect 467925 347520 467930 347576
rect 467986 347520 468340 347576
rect 467925 347518 468340 347520
rect 388529 347515 388595 347518
rect 467925 347515 467991 347518
rect 468334 347516 468340 347518
rect 468404 347516 468410 347580
rect 468526 347578 468586 347654
rect 468661 347712 468708 347716
rect 468772 347714 468778 347716
rect 468661 347656 468666 347712
rect 468661 347652 468708 347656
rect 468772 347654 468818 347714
rect 469765 347712 469812 347716
rect 469876 347714 469882 347716
rect 469765 347656 469770 347712
rect 468772 347652 468778 347654
rect 469765 347652 469812 347656
rect 469876 347654 469922 347714
rect 471237 347712 471284 347716
rect 471348 347714 471354 347716
rect 472065 347714 472131 347717
rect 473353 347716 473419 347717
rect 472198 347714 472204 347716
rect 471237 347656 471242 347712
rect 469876 347652 469882 347654
rect 471237 347652 471284 347656
rect 471348 347654 471394 347714
rect 472065 347712 472204 347714
rect 472065 347656 472070 347712
rect 472126 347656 472204 347712
rect 472065 347654 472204 347656
rect 471348 347652 471354 347654
rect 468661 347651 468727 347652
rect 469765 347651 469831 347652
rect 471237 347651 471303 347652
rect 472065 347651 472131 347654
rect 472198 347652 472204 347654
rect 472268 347652 472274 347716
rect 473302 347714 473308 347716
rect 473262 347654 473308 347714
rect 473372 347712 473419 347716
rect 473414 347656 473419 347712
rect 473302 347652 473308 347654
rect 473372 347652 473419 347656
rect 473353 347651 473419 347652
rect 474365 347716 474431 347717
rect 475653 347716 475719 347717
rect 476941 347716 477007 347717
rect 478045 347716 478111 347717
rect 479149 347716 479215 347717
rect 513373 347716 513439 347717
rect 518341 347716 518407 347717
rect 525885 347716 525951 347717
rect 474365 347712 474412 347716
rect 474476 347714 474482 347716
rect 474365 347656 474370 347712
rect 474365 347652 474412 347656
rect 474476 347654 474522 347714
rect 475653 347712 475700 347716
rect 475764 347714 475770 347716
rect 475653 347656 475658 347712
rect 474476 347652 474482 347654
rect 475653 347652 475700 347656
rect 475764 347654 475810 347714
rect 476941 347712 476988 347716
rect 477052 347714 477058 347716
rect 476941 347656 476946 347712
rect 475764 347652 475770 347654
rect 476941 347652 476988 347656
rect 477052 347654 477098 347714
rect 478045 347712 478092 347716
rect 478156 347714 478162 347716
rect 478045 347656 478050 347712
rect 477052 347652 477058 347654
rect 478045 347652 478092 347656
rect 478156 347654 478202 347714
rect 479149 347712 479196 347716
rect 479260 347714 479266 347716
rect 479149 347656 479154 347712
rect 478156 347652 478162 347654
rect 479149 347652 479196 347656
rect 479260 347654 479306 347714
rect 513373 347712 513420 347716
rect 513484 347714 513490 347716
rect 513373 347656 513378 347712
rect 479260 347652 479266 347654
rect 513373 347652 513420 347656
rect 513484 347654 513530 347714
rect 518341 347712 518388 347716
rect 518452 347714 518458 347716
rect 518341 347656 518346 347712
rect 513484 347652 513490 347654
rect 518341 347652 518388 347656
rect 518452 347654 518498 347714
rect 525885 347712 525932 347716
rect 525996 347714 526002 347716
rect 525885 347656 525890 347712
rect 518452 347652 518458 347654
rect 525885 347652 525932 347656
rect 525996 347654 526042 347714
rect 525996 347652 526002 347654
rect 474365 347651 474431 347652
rect 475653 347651 475719 347652
rect 476941 347651 477007 347652
rect 478045 347651 478111 347652
rect 479149 347651 479215 347652
rect 513373 347651 513439 347652
rect 518341 347651 518407 347652
rect 525885 347651 525951 347652
rect 470358 347578 470364 347580
rect 468526 347518 470364 347578
rect 470358 347516 470364 347518
rect 470428 347516 470434 347580
rect 55806 347380 55812 347444
rect 55876 347442 55882 347444
rect 56593 347442 56659 347445
rect 55876 347440 56659 347442
rect 55876 347384 56598 347440
rect 56654 347384 56659 347440
rect 55876 347382 56659 347384
rect 55876 347380 55882 347382
rect 56593 347379 56659 347382
rect 58198 347380 58204 347444
rect 58268 347442 58274 347444
rect 59353 347442 59419 347445
rect 58268 347440 59419 347442
rect 58268 347384 59358 347440
rect 59414 347384 59419 347440
rect 58268 347382 59419 347384
rect 58268 347380 58274 347382
rect 59353 347379 59419 347382
rect 59486 347380 59492 347444
rect 59556 347442 59562 347444
rect 60825 347442 60891 347445
rect 59556 347440 60891 347442
rect 59556 347384 60830 347440
rect 60886 347384 60891 347440
rect 59556 347382 60891 347384
rect 59556 347380 59562 347382
rect 60825 347379 60891 347382
rect 70894 347380 70900 347444
rect 70964 347442 70970 347444
rect 190637 347442 190703 347445
rect 70964 347440 190703 347442
rect 70964 347384 190642 347440
rect 190698 347384 190703 347440
rect 70964 347382 190703 347384
rect 70964 347380 70970 347382
rect 190637 347379 190703 347382
rect 190821 347442 190887 347445
rect 191557 347442 191623 347445
rect 190821 347440 191623 347442
rect 190821 347384 190826 347440
rect 190882 347384 191562 347440
rect 191618 347384 191623 347440
rect 190821 347382 191623 347384
rect 190821 347379 190887 347382
rect 191557 347379 191623 347382
rect 406193 347442 406259 347445
rect 473486 347442 473492 347444
rect 406193 347440 473492 347442
rect 406193 347384 406198 347440
rect 406254 347384 473492 347440
rect 406193 347382 473492 347384
rect 406193 347379 406259 347382
rect 473486 347380 473492 347382
rect 473556 347380 473562 347444
rect 37181 347308 37247 347309
rect 37181 347306 37228 347308
rect 37100 347304 37228 347306
rect 37292 347306 37298 347308
rect 191465 347306 191531 347309
rect 37292 347304 191531 347306
rect 37100 347248 37186 347304
rect 37292 347248 191470 347304
rect 191526 347248 191531 347304
rect 37100 347246 37228 347248
rect 37181 347244 37228 347246
rect 37292 347246 191531 347248
rect 37292 347244 37298 347246
rect 37181 347243 37247 347244
rect 191465 347243 191531 347246
rect 419625 347306 419691 347309
rect 476062 347306 476068 347308
rect 419625 347304 476068 347306
rect 419625 347248 419630 347304
rect 419686 347248 476068 347304
rect 419625 347246 476068 347248
rect 419625 347243 419691 347246
rect 476062 347244 476068 347246
rect 476132 347244 476138 347308
rect 57094 347108 57100 347172
rect 57164 347170 57170 347172
rect 57973 347170 58039 347173
rect 57164 347168 58039 347170
rect 57164 347112 57978 347168
rect 58034 347112 58039 347168
rect 57164 347110 58039 347112
rect 57164 347108 57170 347110
rect 57973 347107 58039 347110
rect 60590 347108 60596 347172
rect 60660 347170 60666 347172
rect 60733 347170 60799 347173
rect 61929 347170 61995 347173
rect 60660 347168 61995 347170
rect 60660 347112 60738 347168
rect 60794 347112 61934 347168
rect 61990 347112 61995 347168
rect 60660 347110 61995 347112
rect 60660 347108 60666 347110
rect 60733 347107 60799 347110
rect 61929 347107 61995 347110
rect 69289 347170 69355 347173
rect 69790 347170 69796 347172
rect 69289 347168 69796 347170
rect 69289 347112 69294 347168
rect 69350 347112 69796 347168
rect 69289 347110 69796 347112
rect 69289 347107 69355 347110
rect 69790 347108 69796 347110
rect 69860 347108 69866 347172
rect 190637 347170 190703 347173
rect 192334 347170 192340 347172
rect 190637 347168 192340 347170
rect 190637 347112 190642 347168
rect 190698 347112 192340 347168
rect 190637 347110 192340 347112
rect 190637 347107 190703 347110
rect 192334 347108 192340 347110
rect 192404 347108 192410 347172
rect 395705 347170 395771 347173
rect 493358 347170 493364 347172
rect 395705 347168 493364 347170
rect 395705 347112 395710 347168
rect 395766 347112 493364 347168
rect 395705 347110 493364 347112
rect 395705 347107 395771 347110
rect 493358 347108 493364 347110
rect 493428 347108 493434 347172
rect 460565 347036 460631 347037
rect 460565 347032 460612 347036
rect 460676 347034 460682 347036
rect 465257 347034 465323 347037
rect 465942 347034 465948 347036
rect 460565 346976 460570 347032
rect 460565 346972 460612 346976
rect 460676 346974 460722 347034
rect 465257 347032 465948 347034
rect 465257 346976 465262 347032
rect 465318 346976 465948 347032
rect 465257 346974 465948 346976
rect 460676 346972 460682 346974
rect 460565 346971 460631 346972
rect 465257 346971 465323 346974
rect 465942 346972 465948 346974
rect 466012 346972 466018 347036
rect 41781 346900 41847 346901
rect 41781 346896 41828 346900
rect 41892 346898 41898 346900
rect 41781 346840 41786 346896
rect 41781 346836 41828 346840
rect 41892 346838 41938 346898
rect 41892 346836 41898 346838
rect 419574 346836 419580 346900
rect 419644 346898 419650 346900
rect 419809 346898 419875 346901
rect 419644 346896 419875 346898
rect 419644 346840 419814 346896
rect 419870 346840 419875 346896
rect 419644 346838 419875 346840
rect 419644 346836 419650 346838
rect 41781 346835 41847 346836
rect 419809 346835 419875 346838
rect 54518 346700 54524 346764
rect 54588 346762 54594 346764
rect 55121 346762 55187 346765
rect 54588 346760 55187 346762
rect 54588 346704 55126 346760
rect 55182 346704 55187 346760
rect 54588 346702 55187 346704
rect 54588 346700 54594 346702
rect 55121 346699 55187 346702
rect 40534 346428 40540 346492
rect 40604 346490 40610 346492
rect 41321 346490 41387 346493
rect 40604 346488 41387 346490
rect 40604 346432 41326 346488
rect 41382 346432 41387 346488
rect 40604 346430 41387 346432
rect 40604 346428 40610 346430
rect 41321 346427 41387 346430
rect 57973 346490 58039 346493
rect 75453 346490 75519 346493
rect 57973 346488 75519 346490
rect 57973 346432 57978 346488
rect 58034 346432 75458 346488
rect 75514 346432 75519 346488
rect 57973 346430 75519 346432
rect 57973 346427 58039 346430
rect 75453 346427 75519 346430
rect 415853 346354 415919 346357
rect 418613 346354 418679 346357
rect 415853 346352 418679 346354
rect 415853 346296 415858 346352
rect 415914 346296 418618 346352
rect 418674 346296 418679 346352
rect 415853 346294 418679 346296
rect 415853 346291 415919 346294
rect 418613 346291 418679 346294
rect 418613 345674 418679 345677
rect 438853 345674 438919 345677
rect 418613 345672 438919 345674
rect 418613 345616 418618 345672
rect 418674 345616 438858 345672
rect 438914 345616 438919 345672
rect 418613 345614 438919 345616
rect 418613 345611 418679 345614
rect 438853 345611 438919 345614
rect -960 345402 480 345492
rect -960 345342 6930 345402
rect -960 345252 480 345342
rect 6870 345130 6930 345342
rect 18638 345204 18644 345268
rect 18708 345266 18714 345268
rect 41781 345266 41847 345269
rect 42701 345266 42767 345269
rect 18708 345264 42767 345266
rect 18708 345208 41786 345264
rect 41842 345208 42706 345264
rect 42762 345208 42767 345264
rect 18708 345206 42767 345208
rect 18708 345204 18714 345206
rect 41781 345203 41847 345206
rect 42701 345203 42767 345206
rect 191833 345130 191899 345133
rect 6870 345128 191899 345130
rect 6870 345072 191838 345128
rect 191894 345072 191899 345128
rect 6870 345070 191899 345072
rect 191833 345067 191899 345070
rect 583520 338452 584960 338692
rect 150985 335476 151051 335477
rect 551001 335476 551067 335477
rect 150934 335474 150940 335476
rect 150894 335414 150940 335474
rect 151004 335472 151051 335476
rect 550950 335474 550956 335476
rect 151046 335416 151051 335472
rect 150934 335412 150940 335414
rect 151004 335412 151051 335416
rect 550910 335414 550956 335474
rect 551020 335472 551067 335476
rect 551062 335416 551067 335472
rect 550950 335412 550956 335414
rect 551020 335412 551067 335416
rect 150985 335411 151051 335412
rect 551001 335411 551067 335412
rect -960 332196 480 332436
rect 158805 329762 158871 329765
rect 156558 329760 158871 329762
rect 156558 329704 158810 329760
rect 158866 329704 158871 329760
rect 156558 329702 158871 329704
rect 156558 329190 156618 329702
rect 158805 329699 158871 329702
rect 558913 329218 558979 329221
rect 556570 329216 558979 329218
rect 556570 329160 558918 329216
rect 558974 329160 558979 329216
rect 556570 329158 558979 329160
rect 558913 329155 558979 329158
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3877 319290 3943 319293
rect -960 319288 3943 319290
rect -960 319232 3882 319288
rect 3938 319232 3943 319288
rect -960 319230 3943 319232
rect -960 319140 480 319230
rect 3877 319227 3943 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3785 306234 3851 306237
rect -960 306232 3851 306234
rect -960 306176 3790 306232
rect 3846 306176 3851 306232
rect -960 306174 3851 306176
rect -960 306084 480 306174
rect 3785 306171 3851 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3693 293178 3759 293181
rect -960 293176 3759 293178
rect -960 293120 3698 293176
rect 3754 293120 3759 293176
rect -960 293118 3759 293120
rect -960 293028 480 293118
rect 3693 293115 3759 293118
rect 17585 286922 17651 286925
rect 19382 286922 20056 286924
rect 17585 286920 20056 286922
rect 17585 286864 17590 286920
rect 17646 286864 20056 286920
rect 417325 286922 417391 286925
rect 419398 286922 420072 286924
rect 417325 286920 420072 286922
rect 417325 286864 417330 286920
rect 417386 286864 420072 286920
rect 17585 286862 19442 286864
rect 417325 286862 419458 286864
rect 17585 286859 17651 286862
rect 417325 286859 417391 286862
rect 19382 285912 20056 285972
rect 417233 285970 417299 285973
rect 419398 285970 420072 285972
rect 417233 285968 420072 285970
rect 417233 285912 417238 285968
rect 417294 285912 420072 285968
rect 17125 285834 17191 285837
rect 17585 285834 17651 285837
rect 17125 285832 17651 285834
rect 17125 285776 17130 285832
rect 17186 285776 17590 285832
rect 17646 285776 17651 285832
rect 17125 285774 17651 285776
rect 17125 285771 17191 285774
rect 17585 285771 17651 285774
rect 17217 285698 17283 285701
rect 17769 285698 17835 285701
rect 19382 285698 19442 285912
rect 417233 285910 419458 285912
rect 417233 285907 417299 285910
rect 17217 285696 19442 285698
rect 17217 285640 17222 285696
rect 17278 285640 17774 285696
rect 17830 285640 19442 285696
rect 17217 285638 19442 285640
rect 417049 285698 417115 285701
rect 417233 285698 417299 285701
rect 417049 285696 417299 285698
rect 417049 285640 417054 285696
rect 417110 285640 417238 285696
rect 417294 285640 417299 285696
rect 417049 285638 417299 285640
rect 17217 285635 17283 285638
rect 17769 285635 17835 285638
rect 417049 285635 417115 285638
rect 417233 285635 417299 285638
rect 583520 285276 584960 285516
rect 16849 283794 16915 283797
rect 17493 283794 17559 283797
rect 19382 283794 20056 283796
rect 16849 283792 20056 283794
rect 16849 283736 16854 283792
rect 16910 283736 17498 283792
rect 17554 283736 20056 283792
rect 417233 283794 417299 283797
rect 417877 283794 417943 283797
rect 419398 283794 420072 283796
rect 417233 283792 420072 283794
rect 417233 283736 417238 283792
rect 417294 283736 417882 283792
rect 417938 283736 420072 283792
rect 16849 283734 19442 283736
rect 417233 283734 419458 283736
rect 16849 283731 16915 283734
rect 17493 283731 17559 283734
rect 417233 283731 417299 283734
rect 417877 283731 417943 283734
rect 17585 282842 17651 282845
rect 19382 282842 20056 282844
rect 17585 282840 20056 282842
rect 17585 282784 17590 282840
rect 17646 282784 20056 282840
rect 417417 282842 417483 282845
rect 419398 282842 420072 282844
rect 417417 282840 420072 282842
rect 417417 282784 417422 282840
rect 417478 282784 420072 282840
rect 17585 282782 19442 282784
rect 417417 282782 419458 282784
rect 17585 282779 17651 282782
rect 417417 282779 417483 282782
rect 16757 281074 16823 281077
rect 17493 281074 17559 281077
rect 19382 281074 20056 281076
rect 16757 281072 20056 281074
rect 16757 281016 16762 281072
rect 16818 281016 17498 281072
rect 17554 281016 20056 281072
rect 416865 281074 416931 281077
rect 417785 281074 417851 281077
rect 419398 281074 420072 281076
rect 416865 281072 420072 281074
rect 416865 281016 416870 281072
rect 416926 281016 417790 281072
rect 417846 281016 420072 281072
rect 16757 281014 19442 281016
rect 416865 281014 419458 281016
rect 16757 281011 16823 281014
rect 17493 281011 17559 281014
rect 416865 281011 416931 281014
rect 417785 281011 417851 281014
rect -960 279972 480 280212
rect 17309 279986 17375 279989
rect 19382 279986 20056 279988
rect 17309 279984 20056 279986
rect 17309 279928 17314 279984
rect 17370 279928 20056 279984
rect 417693 279986 417759 279989
rect 419398 279986 420072 279988
rect 417693 279984 420072 279986
rect 417693 279928 417698 279984
rect 417754 279928 420072 279984
rect 17309 279926 19442 279928
rect 417693 279926 419458 279928
rect 17309 279923 17375 279926
rect 417693 279923 417759 279926
rect 17401 278762 17467 278765
rect 17677 278762 17743 278765
rect 17401 278760 17743 278762
rect 17401 278704 17406 278760
rect 17462 278704 17682 278760
rect 17738 278704 17743 278760
rect 17401 278702 17743 278704
rect 17401 278699 17467 278702
rect 17677 278699 17743 278702
rect 417601 278762 417667 278765
rect 417734 278762 417740 278764
rect 417601 278760 417740 278762
rect 417601 278704 417606 278760
rect 417662 278704 417740 278760
rect 417601 278702 417740 278704
rect 417601 278699 417667 278702
rect 417734 278700 417740 278702
rect 417804 278700 417810 278764
rect 17677 278218 17743 278221
rect 19382 278218 20056 278220
rect 17677 278216 20056 278218
rect 17677 278160 17682 278216
rect 17738 278160 20056 278216
rect 17677 278158 19442 278160
rect 17677 278155 17743 278158
rect 417734 278156 417740 278220
rect 417804 278218 417810 278220
rect 419398 278218 420072 278220
rect 417804 278160 420072 278218
rect 417804 278158 419458 278160
rect 417804 278156 417810 278158
rect 580809 272234 580875 272237
rect 583520 272234 584960 272324
rect 580809 272232 584960 272234
rect 580809 272176 580814 272232
rect 580870 272176 584960 272232
rect 580809 272174 584960 272176
rect 580809 272171 580875 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3601 267202 3667 267205
rect -960 267200 3667 267202
rect -960 267144 3606 267200
rect 3662 267144 3667 267200
rect -960 267142 3667 267144
rect -960 267052 480 267142
rect 3601 267139 3667 267142
rect 16941 260810 17007 260813
rect 17401 260810 17467 260813
rect 16941 260808 17467 260810
rect 16941 260752 16946 260808
rect 17002 260752 17406 260808
rect 17462 260752 17467 260808
rect 16941 260750 17467 260752
rect 16941 260747 17007 260750
rect 17401 260747 17467 260750
rect 417550 260748 417556 260812
rect 417620 260810 417626 260812
rect 417918 260810 417924 260812
rect 417620 260750 417924 260810
rect 417620 260748 417626 260750
rect 417918 260748 417924 260750
rect 417988 260748 417994 260812
rect 17401 259994 17467 259997
rect 19382 259994 20056 259996
rect 17401 259992 20056 259994
rect 17401 259936 17406 259992
rect 17462 259936 20056 259992
rect 17401 259934 19442 259936
rect 17401 259931 17467 259934
rect 417550 259932 417556 259996
rect 417620 259994 417626 259996
rect 419398 259994 420072 259996
rect 417620 259936 420072 259994
rect 417620 259934 419458 259936
rect 417620 259932 417626 259934
rect 580625 258906 580691 258909
rect 583520 258906 584960 258996
rect 580625 258904 584960 258906
rect 580625 258848 580630 258904
rect 580686 258848 584960 258904
rect 580625 258846 584960 258848
rect 580625 258843 580691 258846
rect 583520 258756 584960 258846
rect 17309 258362 17375 258365
rect 19382 258362 20056 258364
rect 17309 258360 20056 258362
rect 17309 258304 17314 258360
rect 17370 258304 20056 258360
rect 418613 258362 418679 258365
rect 419398 258362 420072 258364
rect 418613 258360 420072 258362
rect 418613 258304 418618 258360
rect 418674 258304 420072 258360
rect 17309 258302 19442 258304
rect 418613 258302 419458 258304
rect 17309 258299 17375 258302
rect 418613 258299 418679 258302
rect 17861 258226 17927 258229
rect 17861 258224 19442 258226
rect 17861 258168 17866 258224
rect 17922 258168 19442 258224
rect 17861 258166 19442 258168
rect 17861 258163 17927 258166
rect 19382 258092 19442 258166
rect 19382 258032 20056 258092
rect 417877 258090 417943 258093
rect 417877 258088 417986 258090
rect 417877 258032 417882 258088
rect 417938 258032 417986 258088
rect 417877 258027 417986 258032
rect 417926 257954 417986 258027
rect 419398 258032 420072 258092
rect 419398 257954 419458 258032
rect 417926 257894 419458 257954
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 191598 250412 191604 250476
rect 191668 250474 191674 250476
rect 308581 250474 308647 250477
rect 191668 250472 308647 250474
rect 191668 250416 308586 250472
rect 308642 250416 308647 250472
rect 191668 250414 308647 250416
rect 191668 250412 191674 250414
rect 308581 250411 308647 250414
rect 18689 249794 18755 249797
rect 93485 249796 93551 249797
rect 18822 249794 18828 249796
rect 18689 249792 18828 249794
rect 18689 249736 18694 249792
rect 18750 249736 18828 249792
rect 18689 249734 18828 249736
rect 18689 249731 18755 249734
rect 18822 249732 18828 249734
rect 18892 249732 18898 249796
rect 93440 249794 93446 249796
rect 93394 249734 93446 249794
rect 93510 249792 93551 249796
rect 93546 249736 93551 249792
rect 93440 249732 93446 249734
rect 93510 249732 93551 249736
rect 93485 249731 93551 249732
rect 95877 249796 95943 249797
rect 98545 249796 98611 249797
rect 103513 249796 103579 249797
rect 105997 249796 106063 249797
rect 108573 249796 108639 249797
rect 111057 249796 111123 249797
rect 95877 249792 95894 249796
rect 95958 249794 95964 249796
rect 98472 249794 98478 249796
rect 95877 249736 95882 249792
rect 95877 249732 95894 249736
rect 95958 249734 96034 249794
rect 98454 249734 98478 249794
rect 95958 249732 95964 249734
rect 98472 249732 98478 249734
rect 98542 249792 98611 249796
rect 98542 249736 98550 249792
rect 98606 249736 98611 249792
rect 98542 249732 98611 249736
rect 103504 249732 103510 249796
rect 103574 249794 103580 249796
rect 105952 249794 105958 249796
rect 103574 249734 103666 249794
rect 105906 249734 105958 249794
rect 106022 249792 106063 249796
rect 108536 249794 108542 249796
rect 106058 249736 106063 249792
rect 103574 249732 103580 249734
rect 105952 249732 105958 249734
rect 106022 249732 106063 249736
rect 108482 249734 108542 249794
rect 108606 249792 108639 249796
rect 110984 249794 110990 249796
rect 108634 249736 108639 249792
rect 108536 249732 108542 249734
rect 108606 249732 108639 249736
rect 110966 249734 110990 249794
rect 110984 249732 110990 249734
rect 111054 249792 111123 249796
rect 111054 249736 111062 249792
rect 111118 249736 111123 249792
rect 111054 249732 111123 249736
rect 95877 249731 95943 249732
rect 98545 249731 98611 249732
rect 103513 249731 103579 249732
rect 105997 249731 106063 249732
rect 108573 249731 108639 249732
rect 111057 249731 111123 249732
rect 405457 249794 405523 249797
rect 485957 249796 486023 249797
rect 488257 249796 488323 249797
rect 491017 249796 491083 249797
rect 495893 249796 495959 249797
rect 498469 249796 498535 249797
rect 500953 249796 501019 249797
rect 503529 249796 503595 249797
rect 468280 249794 468286 249796
rect 405457 249792 468286 249794
rect 405457 249736 405462 249792
rect 405518 249736 468286 249792
rect 405457 249734 468286 249736
rect 405457 249731 405523 249734
rect 468280 249732 468286 249734
rect 468350 249732 468356 249796
rect 485957 249792 485966 249796
rect 486030 249794 486036 249796
rect 485957 249736 485962 249792
rect 485957 249732 485966 249736
rect 486030 249734 486114 249794
rect 488257 249792 488278 249796
rect 488342 249794 488348 249796
rect 490992 249794 490998 249796
rect 488257 249736 488262 249792
rect 486030 249732 486036 249734
rect 488257 249732 488278 249736
rect 488342 249734 488414 249794
rect 490926 249734 490998 249794
rect 491062 249792 491083 249796
rect 495888 249794 495894 249796
rect 491078 249736 491083 249792
rect 488342 249732 488348 249734
rect 490992 249732 490998 249734
rect 491062 249732 491083 249736
rect 495802 249734 495894 249794
rect 495888 249732 495894 249734
rect 495958 249732 495964 249796
rect 498469 249792 498478 249796
rect 498542 249794 498548 249796
rect 500920 249794 500926 249796
rect 498469 249736 498474 249792
rect 498469 249732 498478 249736
rect 498542 249734 498626 249794
rect 500862 249734 500926 249794
rect 500990 249792 501019 249796
rect 503504 249794 503510 249796
rect 501014 249736 501019 249792
rect 498542 249732 498548 249734
rect 500920 249732 500926 249734
rect 500990 249732 501019 249736
rect 503438 249734 503510 249794
rect 503574 249792 503595 249796
rect 503590 249736 503595 249792
rect 503504 249732 503510 249734
rect 503574 249732 503595 249736
rect 485957 249731 486023 249732
rect 488257 249731 488323 249732
rect 491017 249731 491083 249732
rect 495893 249731 495959 249732
rect 498469 249731 498535 249732
rect 500953 249731 501019 249732
rect 503529 249731 503595 249732
rect 50797 249660 50863 249661
rect 53649 249660 53715 249661
rect 56041 249660 56107 249661
rect 58525 249660 58591 249661
rect 113449 249660 113515 249661
rect 50736 249658 50742 249660
rect 50706 249598 50742 249658
rect 50806 249656 50863 249660
rect 53592 249658 53598 249660
rect 50858 249600 50863 249656
rect 50736 249596 50742 249598
rect 50806 249596 50863 249600
rect 53558 249598 53598 249658
rect 53662 249656 53715 249660
rect 53710 249600 53715 249656
rect 53592 249596 53598 249598
rect 53662 249596 53715 249600
rect 56040 249596 56046 249660
rect 56110 249658 56116 249660
rect 58488 249658 58494 249660
rect 56110 249598 56198 249658
rect 58434 249598 58494 249658
rect 58558 249656 58591 249660
rect 113432 249658 113438 249660
rect 58586 249600 58591 249656
rect 56110 249596 56116 249598
rect 58488 249596 58494 249598
rect 58558 249596 58591 249600
rect 113358 249598 113438 249658
rect 113502 249656 113515 249660
rect 113510 249600 113515 249656
rect 113432 249596 113438 249598
rect 113502 249596 113515 249600
rect 50797 249595 50863 249596
rect 53649 249595 53715 249596
rect 56041 249595 56107 249596
rect 58525 249595 58591 249596
rect 113449 249595 113515 249596
rect 115841 249660 115907 249661
rect 120901 249660 120967 249661
rect 115841 249656 115886 249660
rect 115950 249658 115956 249660
rect 115841 249600 115846 249656
rect 115841 249596 115886 249600
rect 115950 249598 115998 249658
rect 120901 249656 120918 249660
rect 120982 249658 120988 249660
rect 402513 249658 402579 249661
rect 470961 249660 471027 249661
rect 483473 249660 483539 249661
rect 505921 249660 505987 249661
rect 508497 249660 508563 249661
rect 515857 249660 515923 249661
rect 520917 249660 520983 249661
rect 461072 249658 461078 249660
rect 120901 249600 120906 249656
rect 115950 249596 115956 249598
rect 120901 249596 120918 249600
rect 120982 249598 121058 249658
rect 402513 249656 461078 249658
rect 402513 249600 402518 249656
rect 402574 249600 461078 249656
rect 402513 249598 461078 249600
rect 120982 249596 120988 249598
rect 115841 249595 115907 249596
rect 120901 249595 120967 249596
rect 402513 249595 402579 249598
rect 461072 249596 461078 249598
rect 461142 249596 461148 249660
rect 470961 249656 471006 249660
rect 471070 249658 471076 249660
rect 470961 249600 470966 249656
rect 470961 249596 471006 249600
rect 471070 249598 471118 249658
rect 483473 249656 483518 249660
rect 483582 249658 483588 249660
rect 483473 249600 483478 249656
rect 471070 249596 471076 249598
rect 483473 249596 483518 249600
rect 483582 249598 483630 249658
rect 505921 249656 505958 249660
rect 506022 249658 506028 249660
rect 505921 249600 505926 249656
rect 483582 249596 483588 249598
rect 505921 249596 505958 249600
rect 506022 249598 506078 249658
rect 508497 249656 508542 249660
rect 508606 249658 508612 249660
rect 508497 249600 508502 249656
rect 506022 249596 506028 249598
rect 508497 249596 508542 249600
rect 508606 249598 508654 249658
rect 515857 249656 515886 249660
rect 515950 249658 515956 249660
rect 520912 249658 520918 249660
rect 515857 249600 515862 249656
rect 508606 249596 508612 249598
rect 515857 249596 515886 249600
rect 515950 249598 516014 249658
rect 520826 249598 520918 249658
rect 515950 249596 515956 249598
rect 520912 249596 520918 249598
rect 520982 249596 520988 249660
rect 470961 249595 471027 249596
rect 483473 249595 483539 249596
rect 505921 249595 505987 249596
rect 508497 249595 508563 249596
rect 515857 249595 515923 249596
rect 520917 249595 520983 249596
rect 418102 249460 418108 249524
rect 418172 249522 418178 249524
rect 418337 249522 418403 249525
rect 418172 249520 418403 249522
rect 418172 249464 418342 249520
rect 418398 249464 418403 249520
rect 418172 249462 418403 249464
rect 418172 249460 418178 249462
rect 418337 249459 418403 249462
rect 418838 249460 418844 249524
rect 418908 249522 418914 249524
rect 476062 249522 476068 249524
rect 418908 249462 476068 249522
rect 418908 249460 418914 249462
rect 476062 249460 476068 249462
rect 476132 249460 476138 249524
rect 473629 249388 473695 249389
rect 473629 249384 473676 249388
rect 473740 249386 473746 249388
rect 473629 249328 473634 249384
rect 473629 249324 473676 249328
rect 473740 249326 473786 249386
rect 473740 249324 473746 249326
rect 473629 249323 473695 249324
rect 35893 248300 35959 248301
rect 35893 248296 35940 248300
rect 36004 248298 36010 248300
rect 36445 248298 36511 248301
rect 37038 248298 37044 248300
rect 35893 248240 35898 248296
rect 35893 248236 35940 248240
rect 36004 248238 36050 248298
rect 36445 248296 37044 248298
rect 36445 248240 36450 248296
rect 36506 248240 37044 248296
rect 36445 248238 37044 248240
rect 36004 248236 36010 248238
rect 35893 248235 35959 248236
rect 36445 248235 36511 248238
rect 37038 248236 37044 248238
rect 37108 248236 37114 248300
rect 38653 248298 38719 248301
rect 44173 248300 44239 248301
rect 46657 248300 46723 248301
rect 50153 248300 50219 248301
rect 61193 248300 61259 248301
rect 39614 248298 39620 248300
rect 38653 248296 39620 248298
rect 38653 248240 38658 248296
rect 38714 248240 39620 248296
rect 38653 248238 39620 248240
rect 38653 248235 38719 248238
rect 39614 248236 39620 248238
rect 39684 248236 39690 248300
rect 44173 248296 44220 248300
rect 44284 248298 44290 248300
rect 46606 248298 46612 248300
rect 44173 248240 44178 248296
rect 44173 248236 44220 248240
rect 44284 248238 44330 248298
rect 46566 248238 46612 248298
rect 46676 248296 46723 248300
rect 50102 248298 50108 248300
rect 46718 248240 46723 248296
rect 44284 248236 44290 248238
rect 46606 248236 46612 248238
rect 46676 248236 46723 248240
rect 50062 248238 50108 248298
rect 50172 248296 50219 248300
rect 61142 248298 61148 248300
rect 50214 248240 50219 248296
rect 50102 248236 50108 248238
rect 50172 248236 50219 248240
rect 61102 248238 61148 248298
rect 61212 248296 61259 248300
rect 61254 248240 61259 248296
rect 61142 248236 61148 248238
rect 61212 248236 61259 248240
rect 44173 248235 44239 248236
rect 46657 248235 46723 248236
rect 50153 248235 50219 248236
rect 61193 248235 61259 248236
rect 61377 248298 61443 248301
rect 61694 248298 61700 248300
rect 61377 248296 61700 248298
rect 61377 248240 61382 248296
rect 61438 248240 61700 248296
rect 61377 248238 61700 248240
rect 61377 248235 61443 248238
rect 61694 248236 61700 248238
rect 61764 248236 61770 248300
rect 62113 248298 62179 248301
rect 63585 248300 63651 248301
rect 62798 248298 62804 248300
rect 62113 248296 62804 248298
rect 62113 248240 62118 248296
rect 62174 248240 62804 248296
rect 62113 248238 62804 248240
rect 62113 248235 62179 248238
rect 62798 248236 62804 248238
rect 62868 248236 62874 248300
rect 63534 248298 63540 248300
rect 63494 248238 63540 248298
rect 63604 248296 63651 248300
rect 63646 248240 63651 248296
rect 63534 248236 63540 248238
rect 63604 248236 63651 248240
rect 63585 248235 63651 248236
rect 64873 248298 64939 248301
rect 65977 248300 66043 248301
rect 65190 248298 65196 248300
rect 64873 248296 65196 248298
rect 64873 248240 64878 248296
rect 64934 248240 65196 248296
rect 64873 248238 65196 248240
rect 64873 248235 64939 248238
rect 65190 248236 65196 248238
rect 65260 248236 65266 248300
rect 65926 248298 65932 248300
rect 65886 248238 65932 248298
rect 65996 248296 66043 248300
rect 66038 248240 66043 248296
rect 65926 248236 65932 248238
rect 65996 248236 66043 248240
rect 65977 248235 66043 248236
rect 67633 248298 67699 248301
rect 70945 248300 71011 248301
rect 68686 248298 68692 248300
rect 67633 248296 68692 248298
rect 67633 248240 67638 248296
rect 67694 248240 68692 248296
rect 67633 248238 68692 248240
rect 67633 248235 67699 248238
rect 68686 248236 68692 248238
rect 68756 248236 68762 248300
rect 70894 248298 70900 248300
rect 70854 248238 70900 248298
rect 70964 248296 71011 248300
rect 71006 248240 71011 248296
rect 70894 248236 70900 248238
rect 70964 248236 71011 248240
rect 73654 248236 73660 248300
rect 73724 248298 73730 248300
rect 73797 248298 73863 248301
rect 73724 248296 73863 248298
rect 73724 248240 73802 248296
rect 73858 248240 73863 248296
rect 73724 248238 73863 248240
rect 73724 248236 73730 248238
rect 70945 248235 71011 248236
rect 73797 248235 73863 248238
rect 77293 248298 77359 248301
rect 78489 248300 78555 248301
rect 83641 248300 83707 248301
rect 78070 248298 78076 248300
rect 77293 248296 78076 248298
rect 77293 248240 77298 248296
rect 77354 248240 78076 248296
rect 77293 248238 78076 248240
rect 77293 248235 77359 248238
rect 78070 248236 78076 248238
rect 78140 248236 78146 248300
rect 78438 248298 78444 248300
rect 78398 248238 78444 248298
rect 78508 248296 78555 248300
rect 83590 248298 83596 248300
rect 78550 248240 78555 248296
rect 78438 248236 78444 248238
rect 78508 248236 78555 248240
rect 83550 248238 83596 248298
rect 83660 248296 83707 248300
rect 83702 248240 83707 248296
rect 83590 248236 83596 248238
rect 83660 248236 83707 248240
rect 125910 248236 125916 248300
rect 125980 248298 125986 248300
rect 389357 248298 389423 248301
rect 443177 248300 443243 248301
rect 443126 248298 443132 248300
rect 125980 248296 389423 248298
rect 125980 248240 389362 248296
rect 389418 248240 389423 248296
rect 125980 248238 389423 248240
rect 443086 248238 443132 248298
rect 443196 248296 443243 248300
rect 443238 248240 443243 248296
rect 125980 248236 125986 248238
rect 78489 248235 78555 248236
rect 83641 248235 83707 248236
rect 389357 248235 389423 248238
rect 443126 248236 443132 248238
rect 443196 248236 443243 248240
rect 443177 248235 443243 248236
rect 447133 248298 447199 248301
rect 448278 248298 448284 248300
rect 447133 248296 448284 248298
rect 447133 248240 447138 248296
rect 447194 248240 448284 248296
rect 447133 248238 448284 248240
rect 447133 248235 447199 248238
rect 448278 248236 448284 248238
rect 448348 248236 448354 248300
rect 448646 248236 448652 248300
rect 448716 248298 448722 248300
rect 449801 248298 449867 248301
rect 450169 248300 450235 248301
rect 450118 248298 450124 248300
rect 448716 248296 449867 248298
rect 448716 248240 449806 248296
rect 449862 248240 449867 248296
rect 448716 248238 449867 248240
rect 450078 248238 450124 248298
rect 450188 248296 450235 248300
rect 450230 248240 450235 248296
rect 448716 248236 448722 248238
rect 449801 248235 449867 248238
rect 450118 248236 450124 248238
rect 450188 248236 450235 248240
rect 450169 248235 450235 248236
rect 450353 248298 450419 248301
rect 450670 248298 450676 248300
rect 450353 248296 450676 248298
rect 450353 248240 450358 248296
rect 450414 248240 450676 248296
rect 450353 248238 450676 248240
rect 450353 248235 450419 248238
rect 450670 248236 450676 248238
rect 450740 248236 450746 248300
rect 451222 248236 451228 248300
rect 451292 248298 451298 248300
rect 451365 248298 451431 248301
rect 451292 248296 451431 248298
rect 451292 248240 451370 248296
rect 451426 248240 451431 248296
rect 451292 248238 451431 248240
rect 451292 248236 451298 248238
rect 451365 248235 451431 248238
rect 452653 248298 452719 248301
rect 453614 248298 453620 248300
rect 452653 248296 453620 248298
rect 452653 248240 452658 248296
rect 452714 248240 453620 248296
rect 452653 248238 453620 248240
rect 452653 248235 452719 248238
rect 453614 248236 453620 248238
rect 453684 248236 453690 248300
rect 455413 248298 455479 248301
rect 456190 248298 456196 248300
rect 455413 248296 456196 248298
rect 455413 248240 455418 248296
rect 455474 248240 456196 248296
rect 455413 248238 456196 248240
rect 455413 248235 455479 248238
rect 456190 248236 456196 248238
rect 456260 248236 456266 248300
rect 462313 248298 462379 248301
rect 462814 248298 462820 248300
rect 462313 248296 462820 248298
rect 462313 248240 462318 248296
rect 462374 248240 462820 248296
rect 462313 248238 462820 248240
rect 462313 248235 462379 248238
rect 462814 248236 462820 248238
rect 462884 248236 462890 248300
rect 467833 248298 467899 248301
rect 468702 248298 468708 248300
rect 467833 248296 468708 248298
rect 467833 248240 467838 248296
rect 467894 248240 468708 248296
rect 467833 248238 468708 248240
rect 467833 248235 467899 248238
rect 468702 248236 468708 248238
rect 468772 248236 468778 248300
rect 37273 248162 37339 248165
rect 38142 248162 38148 248164
rect 37273 248160 38148 248162
rect 37273 248104 37278 248160
rect 37334 248104 38148 248160
rect 37273 248102 38148 248104
rect 37273 248099 37339 248102
rect 38142 248100 38148 248102
rect 38212 248100 38218 248164
rect 40033 248162 40099 248165
rect 40534 248162 40540 248164
rect 40033 248160 40540 248162
rect 40033 248104 40038 248160
rect 40094 248104 40540 248160
rect 40033 248102 40540 248104
rect 40033 248099 40099 248102
rect 40534 248100 40540 248102
rect 40604 248100 40610 248164
rect 41413 248162 41479 248165
rect 43069 248164 43135 248165
rect 45277 248164 45343 248165
rect 47577 248164 47643 248165
rect 41638 248162 41644 248164
rect 41413 248160 41644 248162
rect 41413 248104 41418 248160
rect 41474 248104 41644 248160
rect 41413 248102 41644 248104
rect 41413 248099 41479 248102
rect 41638 248100 41644 248102
rect 41708 248100 41714 248164
rect 43069 248160 43116 248164
rect 43180 248162 43186 248164
rect 43069 248104 43074 248160
rect 43069 248100 43116 248104
rect 43180 248102 43226 248162
rect 45277 248160 45324 248164
rect 45388 248162 45394 248164
rect 47526 248162 47532 248164
rect 45277 248104 45282 248160
rect 43180 248100 43186 248102
rect 45277 248100 45324 248104
rect 45388 248102 45434 248162
rect 47486 248102 47532 248162
rect 47596 248160 47643 248164
rect 47638 248104 47643 248160
rect 45388 248100 45394 248102
rect 47526 248100 47532 248102
rect 47596 248100 47643 248104
rect 48446 248100 48452 248164
rect 48516 248162 48522 248164
rect 180701 248162 180767 248165
rect 48516 248160 180767 248162
rect 48516 248104 180706 248160
rect 180762 248104 180767 248160
rect 48516 248102 180767 248104
rect 48516 248100 48522 248102
rect 43069 248099 43135 248100
rect 45277 248099 45343 248100
rect 47577 248099 47643 248100
rect 180701 248099 180767 248102
rect 403985 248162 404051 248165
rect 478454 248162 478460 248164
rect 403985 248160 478460 248162
rect 403985 248104 403990 248160
rect 404046 248104 478460 248160
rect 403985 248102 478460 248104
rect 403985 248099 404051 248102
rect 478454 248100 478460 248102
rect 478524 248100 478530 248164
rect 19609 248026 19675 248029
rect 60590 248026 60596 248028
rect 19609 248024 60596 248026
rect 19609 247968 19614 248024
rect 19670 247968 60596 248024
rect 19609 247966 60596 247968
rect 19609 247963 19675 247966
rect 60590 247964 60596 247966
rect 60660 247964 60666 248028
rect 63493 248026 63559 248029
rect 81065 248028 81131 248029
rect 86033 248028 86099 248029
rect 88241 248028 88307 248029
rect 91001 248028 91067 248029
rect 63902 248026 63908 248028
rect 63493 248024 63908 248026
rect 63493 247968 63498 248024
rect 63554 247968 63908 248024
rect 63493 247966 63908 247968
rect 48681 247892 48747 247893
rect 58065 247892 58131 247893
rect 48630 247890 48636 247892
rect 48590 247830 48636 247890
rect 48700 247888 48747 247892
rect 58014 247890 58020 247892
rect 48742 247832 48747 247888
rect 48630 247828 48636 247830
rect 48700 247828 48747 247832
rect 57974 247830 58020 247890
rect 58084 247888 58131 247892
rect 58126 247832 58131 247888
rect 58014 247828 58020 247830
rect 58084 247828 58131 247832
rect 48681 247827 48747 247828
rect 58065 247827 58131 247828
rect 59445 247892 59511 247893
rect 59445 247888 59492 247892
rect 59556 247890 59562 247892
rect 60598 247890 60658 247964
rect 63493 247963 63559 247966
rect 63902 247964 63908 247966
rect 63972 247964 63978 248028
rect 79174 248026 79180 248028
rect 64830 247966 79180 248026
rect 64830 247890 64890 247966
rect 79174 247964 79180 247966
rect 79244 247964 79250 248028
rect 81014 248026 81020 248028
rect 80974 247966 81020 248026
rect 81084 248024 81131 248028
rect 85982 248026 85988 248028
rect 81126 247968 81131 248024
rect 81014 247964 81020 247966
rect 81084 247964 81131 247968
rect 85942 247966 85988 248026
rect 86052 248024 86099 248028
rect 88190 248026 88196 248028
rect 86094 247968 86099 248024
rect 85982 247964 85988 247966
rect 86052 247964 86099 247968
rect 88150 247966 88196 248026
rect 88260 248024 88307 248028
rect 90950 248026 90956 248028
rect 88302 247968 88307 248024
rect 88190 247964 88196 247966
rect 88260 247964 88307 247968
rect 90910 247966 90956 248026
rect 91020 248024 91067 248028
rect 91062 247968 91067 248024
rect 90950 247964 90956 247966
rect 91020 247964 91067 247968
rect 100886 247964 100892 248028
rect 100956 248026 100962 248028
rect 101213 248026 101279 248029
rect 100956 248024 101279 248026
rect 100956 247968 101218 248024
rect 101274 247968 101279 248024
rect 100956 247966 101279 247968
rect 100956 247964 100962 247966
rect 81065 247963 81131 247964
rect 86033 247963 86099 247964
rect 88241 247963 88307 247964
rect 91001 247963 91067 247964
rect 101213 247963 101279 247966
rect 118550 247964 118556 248028
rect 118620 248026 118626 248028
rect 174537 248026 174603 248029
rect 118620 248024 174603 248026
rect 118620 247968 174542 248024
rect 174598 247968 174603 248024
rect 118620 247966 174603 247968
rect 118620 247964 118626 247966
rect 174537 247963 174603 247966
rect 402421 248026 402487 248029
rect 460933 248026 460999 248029
rect 402421 248024 460999 248026
rect 402421 247968 402426 248024
rect 402482 247968 460938 248024
rect 460994 247968 460999 248024
rect 402421 247966 460999 247968
rect 402421 247963 402487 247966
rect 460933 247963 460999 247966
rect 461117 248026 461183 248029
rect 461710 248026 461716 248028
rect 461117 248024 461716 248026
rect 461117 247968 461122 248024
rect 461178 247968 461716 248024
rect 461117 247966 461716 247968
rect 461117 247963 461183 247966
rect 461710 247964 461716 247966
rect 461780 247964 461786 248028
rect 465073 248026 465139 248029
rect 465206 248026 465212 248028
rect 465073 248024 465212 248026
rect 465073 247968 465078 248024
rect 465134 247968 465212 248024
rect 465073 247966 465212 247968
rect 465073 247963 465139 247966
rect 465206 247964 465212 247966
rect 465276 247964 465282 248028
rect 66253 247892 66319 247893
rect 67725 247892 67791 247893
rect 68369 247892 68435 247893
rect 76097 247892 76163 247893
rect 66253 247890 66300 247892
rect 59445 247832 59450 247888
rect 59445 247828 59492 247832
rect 59556 247830 59602 247890
rect 60598 247830 64890 247890
rect 66208 247888 66300 247890
rect 66208 247832 66258 247888
rect 66208 247830 66300 247832
rect 59556 247828 59562 247830
rect 66253 247828 66300 247830
rect 66364 247828 66370 247892
rect 67725 247890 67772 247892
rect 67680 247888 67772 247890
rect 67680 247832 67730 247888
rect 67680 247830 67772 247832
rect 67725 247828 67772 247830
rect 67836 247828 67842 247892
rect 68318 247890 68324 247892
rect 68278 247830 68324 247890
rect 68388 247888 68435 247892
rect 76046 247890 76052 247892
rect 68430 247832 68435 247888
rect 68318 247828 68324 247830
rect 68388 247828 68435 247832
rect 76006 247830 76052 247890
rect 76116 247888 76163 247892
rect 76158 247832 76163 247888
rect 76046 247828 76052 247830
rect 76116 247828 76163 247832
rect 123334 247828 123340 247892
rect 123404 247890 123410 247892
rect 171777 247890 171843 247893
rect 123404 247888 171843 247890
rect 123404 247832 171782 247888
rect 171838 247832 171843 247888
rect 123404 247830 171843 247832
rect 123404 247828 123410 247830
rect 59445 247827 59511 247828
rect 66253 247827 66319 247828
rect 67725 247827 67791 247828
rect 68369 247827 68435 247828
rect 76097 247827 76163 247828
rect 171777 247827 171843 247830
rect 405273 247890 405339 247893
rect 461117 247890 461183 247893
rect 463550 247890 463556 247892
rect 405273 247888 461042 247890
rect 405273 247832 405278 247888
rect 405334 247832 461042 247888
rect 405273 247830 461042 247832
rect 405273 247827 405339 247830
rect 18822 247692 18828 247756
rect 18892 247754 18898 247756
rect 29545 247754 29611 247757
rect 18892 247752 29611 247754
rect 18892 247696 29550 247752
rect 29606 247696 29611 247752
rect 18892 247694 29611 247696
rect 18892 247692 18898 247694
rect 29545 247691 29611 247694
rect 74993 247754 75059 247757
rect 75678 247754 75684 247756
rect 74993 247752 75684 247754
rect 74993 247696 74998 247752
rect 75054 247696 75684 247752
rect 74993 247694 75684 247696
rect 74993 247691 75059 247694
rect 75678 247692 75684 247694
rect 75748 247692 75754 247756
rect 75913 247754 75979 247757
rect 76966 247754 76972 247756
rect 75913 247752 76972 247754
rect 75913 247696 75918 247752
rect 75974 247696 76972 247752
rect 75913 247694 76972 247696
rect 75913 247691 75979 247694
rect 76966 247692 76972 247694
rect 77036 247692 77042 247756
rect 402605 247754 402671 247757
rect 458398 247754 458404 247756
rect 402605 247752 458404 247754
rect 402605 247696 402610 247752
rect 402666 247696 458404 247752
rect 402605 247694 458404 247696
rect 402605 247691 402671 247694
rect 458398 247692 458404 247694
rect 458468 247692 458474 247756
rect 460982 247754 461042 247830
rect 461117 247888 463556 247890
rect 461117 247832 461122 247888
rect 461178 247832 463556 247888
rect 461117 247830 463556 247832
rect 461117 247827 461183 247830
rect 463550 247828 463556 247830
rect 463620 247828 463626 247892
rect 463693 247890 463759 247893
rect 463918 247890 463924 247892
rect 463693 247888 463924 247890
rect 463693 247832 463698 247888
rect 463754 247832 463924 247888
rect 463693 247830 463924 247832
rect 463693 247827 463759 247830
rect 463918 247828 463924 247830
rect 463988 247828 463994 247892
rect 469213 247890 469279 247893
rect 469806 247890 469812 247892
rect 469213 247888 469812 247890
rect 469213 247832 469218 247888
rect 469274 247832 469812 247888
rect 469213 247830 469812 247832
rect 469213 247827 469279 247830
rect 469806 247828 469812 247830
rect 469876 247828 469882 247892
rect 473353 247890 473419 247893
rect 474406 247890 474412 247892
rect 473353 247888 474412 247890
rect 473353 247832 473358 247888
rect 473414 247832 474412 247888
rect 473353 247830 474412 247832
rect 473353 247827 473419 247830
rect 474406 247828 474412 247830
rect 474476 247828 474482 247892
rect 465942 247754 465948 247756
rect 460982 247694 465948 247754
rect 465942 247692 465948 247694
rect 466012 247692 466018 247756
rect 466453 247754 466519 247757
rect 467598 247754 467604 247756
rect 466453 247752 467604 247754
rect 466453 247696 466458 247752
rect 466514 247696 467604 247752
rect 466453 247694 467604 247696
rect 466453 247691 466519 247694
rect 467598 247692 467604 247694
rect 467668 247692 467674 247756
rect 478873 247754 478939 247757
rect 479190 247754 479196 247756
rect 478873 247752 479196 247754
rect 478873 247696 478878 247752
rect 478934 247696 479196 247752
rect 478873 247694 479196 247696
rect 478873 247691 478939 247694
rect 479190 247692 479196 247694
rect 479260 247692 479266 247756
rect 18638 247556 18644 247620
rect 18708 247618 18714 247620
rect 38101 247618 38167 247621
rect 18708 247616 38167 247618
rect 18708 247560 38106 247616
rect 38162 247560 38167 247616
rect 18708 247558 38167 247560
rect 18708 247556 18714 247558
rect 38101 247555 38167 247558
rect 71773 247618 71839 247621
rect 72182 247618 72188 247620
rect 71773 247616 72188 247618
rect 71773 247560 71778 247616
rect 71834 247560 72188 247616
rect 71773 247558 72188 247560
rect 71773 247555 71839 247558
rect 72182 247556 72188 247558
rect 72252 247556 72258 247620
rect 414473 247618 414539 247621
rect 417785 247618 417851 247621
rect 455873 247620 455939 247621
rect 455822 247618 455828 247620
rect 414473 247616 451290 247618
rect 414473 247560 414478 247616
rect 414534 247560 417790 247616
rect 417846 247560 451290 247616
rect 414473 247558 451290 247560
rect 455782 247558 455828 247618
rect 455892 247616 455939 247620
rect 460606 247618 460612 247620
rect 455934 247560 455939 247616
rect 414473 247555 414539 247558
rect 417785 247555 417851 247558
rect 51390 247420 51396 247484
rect 51460 247482 51466 247484
rect 52361 247482 52427 247485
rect 51460 247480 52427 247482
rect 51460 247424 52366 247480
rect 52422 247424 52427 247480
rect 51460 247422 52427 247424
rect 51460 247420 51466 247422
rect 52361 247419 52427 247422
rect 69013 247482 69079 247485
rect 69790 247482 69796 247484
rect 69013 247480 69796 247482
rect 69013 247424 69018 247480
rect 69074 247424 69796 247480
rect 69013 247422 69796 247424
rect 69013 247419 69079 247422
rect 69790 247420 69796 247422
rect 69860 247420 69866 247484
rect 451230 247482 451290 247558
rect 455822 247556 455828 247558
rect 455892 247556 455939 247560
rect 455873 247555 455939 247556
rect 457670 247558 460612 247618
rect 457670 247482 457730 247558
rect 460606 247556 460612 247558
rect 460676 247618 460682 247620
rect 462221 247618 462287 247621
rect 460676 247616 462287 247618
rect 460676 247560 462226 247616
rect 462282 247560 462287 247616
rect 460676 247558 462287 247560
rect 460676 247556 460682 247558
rect 462221 247555 462287 247558
rect 465073 247618 465139 247621
rect 466310 247618 466316 247620
rect 465073 247616 466316 247618
rect 465073 247560 465078 247616
rect 465134 247560 466316 247616
rect 465073 247558 466316 247560
rect 465073 247555 465139 247558
rect 466310 247556 466316 247558
rect 466380 247556 466386 247620
rect 470777 247618 470843 247621
rect 471278 247618 471284 247620
rect 470777 247616 471284 247618
rect 470777 247560 470782 247616
rect 470838 247560 471284 247616
rect 470777 247558 471284 247560
rect 470777 247555 470843 247558
rect 471278 247556 471284 247558
rect 471348 247556 471354 247620
rect 457989 247482 458055 247485
rect 475694 247482 475700 247484
rect 451230 247422 457730 247482
rect 457854 247480 475700 247482
rect 457854 247424 457994 247480
rect 458050 247424 475700 247480
rect 457854 247422 475700 247424
rect 53414 247284 53420 247348
rect 53484 247346 53490 247348
rect 53741 247346 53807 247349
rect 53484 247344 53807 247346
rect 53484 247288 53746 247344
rect 53802 247288 53807 247344
rect 53484 247286 53807 247288
rect 53484 247284 53490 247286
rect 53741 247283 53807 247286
rect 70393 247346 70459 247349
rect 71262 247346 71268 247348
rect 70393 247344 71268 247346
rect 70393 247288 70398 247344
rect 70454 247288 71268 247344
rect 70393 247286 71268 247288
rect 70393 247283 70459 247286
rect 71262 247284 71268 247286
rect 71332 247284 71338 247348
rect 73245 247346 73311 247349
rect 74390 247346 74396 247348
rect 73245 247344 74396 247346
rect 73245 247288 73250 247344
rect 73306 247288 74396 247344
rect 73245 247286 74396 247288
rect 73245 247283 73311 247286
rect 74390 247284 74396 247286
rect 74460 247284 74466 247348
rect 436093 247346 436159 247349
rect 437054 247346 437060 247348
rect 436093 247344 437060 247346
rect 436093 247288 436098 247344
rect 436154 247288 437060 247344
rect 436093 247286 437060 247288
rect 436093 247283 436159 247286
rect 437054 247284 437060 247286
rect 437124 247284 437130 247348
rect 457110 247284 457116 247348
rect 457180 247346 457186 247348
rect 457854 247346 457914 247422
rect 457989 247419 458055 247422
rect 475694 247420 475700 247422
rect 475764 247420 475770 247484
rect 476113 247482 476179 247485
rect 476982 247482 476988 247484
rect 476113 247480 476988 247482
rect 476113 247424 476118 247480
rect 476174 247424 476988 247480
rect 476113 247422 476988 247424
rect 476113 247419 476179 247422
rect 476982 247420 476988 247422
rect 477052 247420 477058 247484
rect 457180 247286 457914 247346
rect 459461 247348 459527 247349
rect 459461 247344 459508 247348
rect 459572 247346 459578 247348
rect 471973 247346 472039 247349
rect 473353 247348 473419 247349
rect 472198 247346 472204 247348
rect 459461 247288 459466 247344
rect 457180 247284 457186 247286
rect 459461 247284 459508 247288
rect 459572 247286 459618 247346
rect 471973 247344 472204 247346
rect 471973 247288 471978 247344
rect 472034 247288 472204 247344
rect 471973 247286 472204 247288
rect 459572 247284 459578 247286
rect 459461 247283 459527 247284
rect 471973 247283 472039 247286
rect 472198 247284 472204 247286
rect 472268 247284 472274 247348
rect 473302 247284 473308 247348
rect 473372 247346 473419 247348
rect 477493 247346 477559 247349
rect 478086 247346 478092 247348
rect 473372 247344 473464 247346
rect 473414 247288 473464 247344
rect 473372 247286 473464 247288
rect 477493 247344 478092 247346
rect 477493 247288 477498 247344
rect 477554 247288 478092 247344
rect 477493 247286 478092 247288
rect 473372 247284 473419 247286
rect 473353 247283 473419 247284
rect 477493 247283 477559 247286
rect 478086 247284 478092 247286
rect 478156 247284 478162 247348
rect 73153 247210 73219 247213
rect 73286 247210 73292 247212
rect 73153 247208 73292 247210
rect 73153 247152 73158 247208
rect 73214 247152 73292 247208
rect 73153 247150 73292 247152
rect 73153 247147 73219 247150
rect 73286 247148 73292 247150
rect 73356 247148 73362 247212
rect 398097 247210 398163 247213
rect 518382 247210 518388 247212
rect 398097 247208 518388 247210
rect 398097 247152 398102 247208
rect 398158 247152 518388 247208
rect 398097 247150 518388 247152
rect 398097 247147 398163 247150
rect 518382 247148 518388 247150
rect 518452 247148 518458 247212
rect 52361 247076 52427 247077
rect 52310 247074 52316 247076
rect 52270 247014 52316 247074
rect 52380 247072 52427 247076
rect 52422 247016 52427 247072
rect 52310 247012 52316 247014
rect 52380 247012 52427 247016
rect 54518 247012 54524 247076
rect 54588 247074 54594 247076
rect 55121 247074 55187 247077
rect 54588 247072 55187 247074
rect 54588 247016 55126 247072
rect 55182 247016 55187 247072
rect 54588 247014 55187 247016
rect 54588 247012 54594 247014
rect 52361 247011 52427 247012
rect 55121 247011 55187 247014
rect 55806 247012 55812 247076
rect 55876 247074 55882 247076
rect 56501 247074 56567 247077
rect 55876 247072 56567 247074
rect 55876 247016 56506 247072
rect 56562 247016 56567 247072
rect 55876 247014 56567 247016
rect 55876 247012 55882 247014
rect 56501 247011 56567 247014
rect 57094 247012 57100 247076
rect 57164 247074 57170 247076
rect 57973 247074 58039 247077
rect 63217 247074 63283 247077
rect 436185 247076 436251 247077
rect 436134 247074 436140 247076
rect 57164 247072 63283 247074
rect 57164 247016 57978 247072
rect 58034 247016 63222 247072
rect 63278 247016 63283 247072
rect 57164 247014 63283 247016
rect 436094 247014 436140 247074
rect 436204 247072 436251 247076
rect 436246 247016 436251 247072
rect 57164 247012 57170 247014
rect 57973 247011 58039 247014
rect 63217 247011 63283 247014
rect 436134 247012 436140 247014
rect 436204 247012 436251 247016
rect 436185 247011 436251 247012
rect 437473 247074 437539 247077
rect 438158 247074 438164 247076
rect 437473 247072 438164 247074
rect 437473 247016 437478 247072
rect 437534 247016 438164 247072
rect 437473 247014 438164 247016
rect 437473 247011 437539 247014
rect 438158 247012 438164 247014
rect 438228 247012 438234 247076
rect 438853 247074 438919 247077
rect 439630 247074 439636 247076
rect 438853 247072 439636 247074
rect 438853 247016 438858 247072
rect 438914 247016 439636 247072
rect 438853 247014 439636 247016
rect 438853 247011 438919 247014
rect 439630 247012 439636 247014
rect 439700 247012 439706 247076
rect 440233 247074 440299 247077
rect 441613 247076 441679 247077
rect 444281 247076 444347 247077
rect 440550 247074 440556 247076
rect 440233 247072 440556 247074
rect 440233 247016 440238 247072
rect 440294 247016 440556 247072
rect 440233 247014 440556 247016
rect 440233 247011 440299 247014
rect 440550 247012 440556 247014
rect 440620 247012 440626 247076
rect 441613 247072 441660 247076
rect 441724 247074 441730 247076
rect 444230 247074 444236 247076
rect 441613 247016 441618 247072
rect 441613 247012 441660 247016
rect 441724 247014 441770 247074
rect 444190 247014 444236 247074
rect 444300 247072 444347 247076
rect 444342 247016 444347 247072
rect 441724 247012 441730 247014
rect 444230 247012 444236 247014
rect 444300 247012 444347 247016
rect 445518 247012 445524 247076
rect 445588 247074 445594 247076
rect 445661 247074 445727 247077
rect 445588 247072 445727 247074
rect 445588 247016 445666 247072
rect 445722 247016 445727 247072
rect 445588 247014 445727 247016
rect 445588 247012 445594 247014
rect 441613 247011 441679 247012
rect 444281 247011 444347 247012
rect 445661 247011 445727 247014
rect 446622 247012 446628 247076
rect 446692 247074 446698 247076
rect 447041 247074 447107 247077
rect 446692 247072 447107 247074
rect 446692 247016 447046 247072
rect 447102 247016 447107 247072
rect 446692 247014 447107 247016
rect 446692 247012 446698 247014
rect 447041 247011 447107 247014
rect 447726 247012 447732 247076
rect 447796 247074 447802 247076
rect 448421 247074 448487 247077
rect 447796 247072 448487 247074
rect 447796 247016 448426 247072
rect 448482 247016 448487 247072
rect 447796 247014 448487 247016
rect 447796 247012 447802 247014
rect 448421 247011 448487 247014
rect 452326 247012 452332 247076
rect 452396 247074 452402 247076
rect 452561 247074 452627 247077
rect 452396 247072 452627 247074
rect 452396 247016 452566 247072
rect 452622 247016 452627 247072
rect 452396 247014 452627 247016
rect 452396 247012 452402 247014
rect 452561 247011 452627 247014
rect 453430 247012 453436 247076
rect 453500 247074 453506 247076
rect 453941 247074 454007 247077
rect 453500 247072 454007 247074
rect 453500 247016 453946 247072
rect 454002 247016 454007 247072
rect 453500 247014 454007 247016
rect 453500 247012 453506 247014
rect 453941 247011 454007 247014
rect 454534 247012 454540 247076
rect 454604 247074 454610 247076
rect 455321 247074 455387 247077
rect 458081 247076 458147 247077
rect 458030 247074 458036 247076
rect 454604 247072 455387 247074
rect 454604 247016 455326 247072
rect 455382 247016 455387 247072
rect 454604 247014 455387 247016
rect 457990 247014 458036 247074
rect 458100 247072 458147 247076
rect 458142 247016 458147 247072
rect 454604 247012 454610 247014
rect 455321 247011 455387 247014
rect 458030 247012 458036 247014
rect 458100 247012 458147 247016
rect 458081 247011 458147 247012
rect 480529 247074 480595 247077
rect 480846 247074 480852 247076
rect 480529 247072 480852 247074
rect 480529 247016 480534 247072
rect 480590 247016 480852 247072
rect 480529 247014 480852 247016
rect 480529 247011 480595 247014
rect 480846 247012 480852 247014
rect 480916 247012 480922 247076
rect 492673 247074 492739 247077
rect 493358 247074 493364 247076
rect 492673 247072 493364 247074
rect 492673 247016 492678 247072
rect 492734 247016 493364 247072
rect 492673 247014 493364 247016
rect 492673 247011 492739 247014
rect 493358 247012 493364 247014
rect 493428 247012 493434 247076
rect 510613 247074 510679 247077
rect 513373 247076 513439 247077
rect 511022 247074 511028 247076
rect 510613 247072 511028 247074
rect 510613 247016 510618 247072
rect 510674 247016 511028 247072
rect 510613 247014 511028 247016
rect 510613 247011 510679 247014
rect 511022 247012 511028 247014
rect 511092 247012 511098 247076
rect 513373 247074 513420 247076
rect 513328 247072 513420 247074
rect 513328 247016 513378 247072
rect 513328 247014 513420 247016
rect 513373 247012 513420 247014
rect 513484 247012 513490 247076
rect 523033 247074 523099 247077
rect 523350 247074 523356 247076
rect 523033 247072 523356 247074
rect 523033 247016 523038 247072
rect 523094 247016 523356 247072
rect 523033 247014 523356 247016
rect 513373 247011 513439 247012
rect 523033 247011 523099 247014
rect 523350 247012 523356 247014
rect 523420 247012 523426 247076
rect 525793 247074 525859 247077
rect 525926 247074 525932 247076
rect 525793 247072 525932 247074
rect 525793 247016 525798 247072
rect 525854 247016 525932 247072
rect 525793 247014 525932 247016
rect 525793 247011 525859 247014
rect 525926 247012 525932 247014
rect 525996 247012 526002 247076
rect 580533 245578 580599 245581
rect 583520 245578 584960 245668
rect 580533 245576 584960 245578
rect 580533 245520 580538 245576
rect 580594 245520 584960 245576
rect 580533 245518 584960 245520
rect 580533 245515 580599 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 419942 238580 419948 238644
rect 420012 238642 420018 238644
rect 459553 238642 459619 238645
rect 420012 238640 459619 238642
rect 420012 238584 459558 238640
rect 459614 238584 459619 238640
rect 420012 238582 459619 238584
rect 420012 238580 420018 238582
rect 459553 238579 459619 238582
rect 418981 235922 419047 235925
rect 419206 235922 419212 235924
rect 418981 235920 419212 235922
rect 418981 235864 418986 235920
rect 419042 235864 419212 235920
rect 418981 235862 419212 235864
rect 418981 235859 419047 235862
rect 419206 235860 419212 235862
rect 419276 235922 419282 235924
rect 441613 235922 441679 235925
rect 419276 235920 441679 235922
rect 419276 235864 441618 235920
rect 441674 235864 441679 235920
rect 419276 235862 441679 235864
rect 419276 235860 419282 235862
rect 441613 235859 441679 235862
rect 419574 235724 419580 235788
rect 419644 235786 419650 235788
rect 440233 235786 440299 235789
rect 419644 235784 440299 235786
rect 419644 235728 440238 235784
rect 440294 235728 440299 235784
rect 419644 235726 440299 235728
rect 419644 235724 419650 235726
rect 440233 235723 440299 235726
rect 419165 235650 419231 235653
rect 438853 235650 438919 235653
rect 419165 235648 438919 235650
rect 419165 235592 419170 235648
rect 419226 235592 438858 235648
rect 438914 235592 438919 235648
rect 419165 235590 438919 235592
rect 419165 235587 419231 235590
rect 438853 235587 438919 235590
rect 418613 235514 418679 235517
rect 437473 235514 437539 235517
rect 418613 235512 437539 235514
rect 418613 235456 418618 235512
rect 418674 235456 437478 235512
rect 437534 235456 437539 235512
rect 418613 235454 437539 235456
rect 418613 235451 418679 235454
rect 437473 235451 437539 235454
rect 550817 235108 550883 235109
rect 550766 235106 550772 235108
rect 550726 235046 550772 235106
rect 550836 235104 550883 235108
rect 550878 235048 550883 235104
rect 550766 235044 550772 235046
rect 550836 235044 550883 235048
rect 550817 235043 550883 235044
rect 150433 234698 150499 234701
rect 150750 234698 150756 234700
rect 150433 234696 150756 234698
rect 150433 234640 150438 234696
rect 150494 234640 150756 234696
rect 150433 234638 150756 234640
rect 150433 234635 150499 234638
rect 150750 234636 150756 234638
rect 150820 234636 150826 234700
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 158713 229258 158779 229261
rect 557625 229258 557691 229261
rect 558913 229258 558979 229261
rect 156558 229256 158779 229258
rect 156558 229200 158718 229256
rect 158774 229200 158779 229256
rect 156558 229198 158779 229200
rect 156558 229190 156618 229198
rect 158713 229195 158779 229198
rect 556570 229256 558979 229258
rect 556570 229200 557630 229256
rect 557686 229200 558918 229256
rect 558974 229200 558979 229256
rect 556570 229198 558979 229200
rect 556570 229190 556630 229198
rect 557625 229195 557691 229198
rect 558913 229195 558979 229198
rect -960 227884 480 228124
rect 579981 219058 580047 219061
rect 583520 219058 584960 219148
rect 579981 219056 584960 219058
rect 579981 219000 579986 219056
rect 580042 219000 584960 219056
rect 579981 218998 584960 219000
rect 579981 218995 580047 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580441 205730 580507 205733
rect 583520 205730 584960 205820
rect 580441 205728 584960 205730
rect 580441 205672 580446 205728
rect 580502 205672 584960 205728
rect 580441 205670 584960 205672
rect 580441 205667 580507 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 16757 186962 16823 186965
rect 17125 186962 17191 186965
rect 417325 186962 417391 186965
rect 417877 186962 417943 186965
rect 16757 186960 19442 186962
rect 16757 186904 16762 186960
rect 16818 186904 17130 186960
rect 17186 186924 19442 186960
rect 417325 186960 419458 186962
rect 17186 186904 20056 186924
rect 16757 186902 20056 186904
rect 16757 186899 16823 186902
rect 17125 186899 17191 186902
rect 19382 186864 20056 186902
rect 417325 186904 417330 186960
rect 417386 186904 417882 186960
rect 417938 186924 419458 186960
rect 417938 186904 420072 186924
rect 417325 186902 420072 186904
rect 417325 186899 417391 186902
rect 417877 186899 417943 186902
rect 419398 186864 420072 186902
rect 17125 186010 17191 186013
rect 17769 186010 17835 186013
rect 417049 186010 417115 186013
rect 17125 186008 19442 186010
rect 17125 185952 17130 186008
rect 17186 185952 17774 186008
rect 17830 185972 19442 186008
rect 417049 186008 419458 186010
rect 17830 185952 20056 185972
rect 17125 185950 20056 185952
rect 17125 185947 17191 185950
rect 17769 185947 17835 185950
rect 19382 185912 20056 185950
rect 417049 185952 417054 186008
rect 417110 185972 419458 186008
rect 417110 185952 420072 185972
rect 417049 185950 420072 185952
rect 417049 185947 417115 185950
rect 419398 185912 420072 185950
rect 16849 183834 16915 183837
rect 417233 183834 417299 183837
rect 417969 183834 418035 183837
rect 16849 183832 19442 183834
rect 16849 183776 16854 183832
rect 16910 183796 19442 183832
rect 417233 183832 419458 183834
rect 16910 183776 20056 183796
rect 16849 183774 20056 183776
rect 16849 183771 16915 183774
rect 19382 183736 20056 183774
rect 417233 183776 417238 183832
rect 417294 183776 417974 183832
rect 418030 183796 419458 183832
rect 418030 183776 420072 183796
rect 417233 183774 420072 183776
rect 417233 183771 417299 183774
rect 417969 183771 418035 183774
rect 419398 183736 420072 183774
rect 17585 182882 17651 182885
rect 417417 182882 417483 182885
rect 17585 182880 19442 182882
rect 17585 182824 17590 182880
rect 17646 182844 19442 182880
rect 417417 182880 419458 182882
rect 17646 182824 20056 182844
rect 17585 182822 20056 182824
rect 17585 182819 17651 182822
rect 19382 182784 20056 182822
rect 417417 182824 417422 182880
rect 417478 182844 419458 182880
rect 417478 182824 420072 182844
rect 417417 182822 420072 182824
rect 417417 182819 417483 182822
rect 419398 182784 420072 182822
rect 416865 182066 416931 182069
rect 417233 182066 417299 182069
rect 416865 182064 417299 182066
rect 416865 182008 416870 182064
rect 416926 182008 417238 182064
rect 417294 182008 417299 182064
rect 416865 182006 417299 182008
rect 416865 182003 416931 182006
rect 417233 182003 417299 182006
rect 17493 181114 17559 181117
rect 417233 181114 417299 181117
rect 17493 181112 19442 181114
rect 17493 181056 17498 181112
rect 17554 181076 19442 181112
rect 417233 181112 419458 181114
rect 17554 181056 20056 181076
rect 17493 181054 20056 181056
rect 17493 181051 17559 181054
rect 19382 181016 20056 181054
rect 417233 181056 417238 181112
rect 417294 181076 419458 181112
rect 417294 181056 420072 181076
rect 417233 181054 420072 181056
rect 417233 181051 417299 181054
rect 419398 181016 420072 181054
rect 17861 180026 17927 180029
rect 417509 180026 417575 180029
rect 17861 180024 19442 180026
rect 17861 179968 17866 180024
rect 17922 179988 19442 180024
rect 417509 180024 419458 180026
rect 17922 179968 20056 179988
rect 17861 179966 20056 179968
rect 17861 179963 17927 179966
rect 19382 179928 20056 179966
rect 417509 179968 417514 180024
rect 417570 179988 419458 180024
rect 417570 179968 420072 179988
rect 417509 179966 420072 179968
rect 417509 179963 417575 179966
rect 419398 179928 420072 179966
rect 17217 179482 17283 179485
rect 17861 179482 17927 179485
rect 17217 179480 17927 179482
rect 17217 179424 17222 179480
rect 17278 179424 17866 179480
rect 17922 179424 17927 179480
rect 17217 179422 17927 179424
rect 17217 179419 17283 179422
rect 17861 179419 17927 179422
rect 417509 179482 417575 179485
rect 417918 179482 417924 179484
rect 417509 179480 417924 179482
rect 417509 179424 417514 179480
rect 417570 179424 417924 179480
rect 417509 179422 417924 179424
rect 417509 179419 417575 179422
rect 417918 179420 417924 179422
rect 417988 179420 417994 179484
rect 580073 179210 580139 179213
rect 583520 179210 584960 179300
rect 580073 179208 584960 179210
rect 580073 179152 580078 179208
rect 580134 179152 584960 179208
rect 580073 179150 584960 179152
rect 580073 179147 580139 179150
rect 583520 179060 584960 179150
rect 17769 178258 17835 178261
rect 17769 178256 19442 178258
rect 17769 178200 17774 178256
rect 17830 178220 19442 178256
rect 17830 178200 20056 178220
rect 17769 178198 20056 178200
rect 17769 178195 17835 178198
rect 19382 178160 20056 178198
rect 417734 178196 417740 178260
rect 417804 178258 417810 178260
rect 417804 178220 419458 178258
rect 417804 178198 420072 178220
rect 417804 178196 417810 178198
rect 419398 178160 420072 178198
rect -960 175796 480 176036
rect 580533 165882 580599 165885
rect 583520 165882 584960 165972
rect 580533 165880 584960 165882
rect 580533 165824 580538 165880
rect 580594 165824 584960 165880
rect 580533 165822 584960 165824
rect 580533 165819 580599 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 17401 160034 17467 160037
rect 17401 160032 19442 160034
rect 17401 159976 17406 160032
rect 17462 159996 19442 160032
rect 17462 159976 20056 159996
rect 17401 159974 20056 159976
rect 17401 159971 17467 159974
rect 19382 159936 20056 159974
rect 417550 159972 417556 160036
rect 417620 160034 417626 160036
rect 417620 159996 419458 160034
rect 417620 159974 420072 159996
rect 417620 159972 417626 159974
rect 419398 159936 420072 159974
rect 17309 158402 17375 158405
rect 417601 158402 417667 158405
rect 17309 158400 19442 158402
rect 17309 158344 17314 158400
rect 17370 158364 19442 158400
rect 417601 158400 419458 158402
rect 17370 158344 20056 158364
rect 17309 158342 20056 158344
rect 17309 158339 17375 158342
rect 19382 158304 20056 158342
rect 417601 158344 417606 158400
rect 417662 158364 419458 158400
rect 417662 158344 420072 158364
rect 417601 158342 420072 158344
rect 417601 158339 417667 158342
rect 419398 158304 420072 158342
rect 19006 158068 19012 158132
rect 19076 158130 19082 158132
rect 417693 158130 417759 158133
rect 19076 158092 19626 158130
rect 417693 158128 419458 158130
rect 19076 158070 20056 158092
rect 19076 158068 19082 158070
rect 19566 158032 20056 158070
rect 417693 158072 417698 158128
rect 417754 158092 419458 158128
rect 417754 158072 420072 158092
rect 417693 158070 420072 158072
rect 417693 158067 417759 158070
rect 419398 158032 420072 158070
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 580349 152627 580415 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 458081 149836 458147 149837
rect 478505 149836 478571 149837
rect 3366 149834 3372 149836
rect -960 149774 3372 149834
rect -960 149684 480 149774
rect 3366 149772 3372 149774
rect 3436 149772 3442 149836
rect 458080 149834 458086 149836
rect 457994 149774 458086 149834
rect 458080 149772 458086 149774
rect 458150 149772 458156 149836
rect 478480 149834 478486 149836
rect 478414 149774 478486 149834
rect 478550 149832 478571 149836
rect 478566 149776 478571 149832
rect 478480 149772 478486 149774
rect 478550 149772 478571 149776
rect 458081 149771 458147 149772
rect 478505 149771 478571 149772
rect 480897 149836 480963 149837
rect 483473 149836 483539 149837
rect 485957 149836 486023 149837
rect 480897 149832 480934 149836
rect 480998 149834 481004 149836
rect 480897 149776 480902 149832
rect 480897 149772 480934 149776
rect 480998 149774 481054 149834
rect 483473 149832 483518 149836
rect 483582 149834 483588 149836
rect 483473 149776 483478 149832
rect 480998 149772 481004 149774
rect 483473 149772 483518 149776
rect 483582 149774 483630 149834
rect 485957 149832 485966 149836
rect 486030 149834 486036 149836
rect 485957 149776 485962 149832
rect 483582 149772 483588 149774
rect 485957 149772 485966 149776
rect 486030 149774 486114 149834
rect 486030 149772 486036 149774
rect 480897 149771 480963 149772
rect 483473 149771 483539 149772
rect 485957 149771 486023 149772
rect 440049 149698 440115 149701
rect 488257 149700 488323 149701
rect 491017 149700 491083 149701
rect 495893 149700 495959 149701
rect 503529 149700 503595 149701
rect 440536 149698 440542 149700
rect 440049 149696 440542 149698
rect 440049 149640 440054 149696
rect 440110 149640 440542 149696
rect 440049 149638 440542 149640
rect 440049 149635 440115 149638
rect 440536 149636 440542 149638
rect 440606 149636 440612 149700
rect 488257 149696 488278 149700
rect 488342 149698 488348 149700
rect 490992 149698 490998 149700
rect 488257 149640 488262 149696
rect 488257 149636 488278 149640
rect 488342 149638 488414 149698
rect 490926 149638 490998 149698
rect 491062 149696 491083 149700
rect 495888 149698 495894 149700
rect 491078 149640 491083 149696
rect 488342 149636 488348 149638
rect 490992 149636 490998 149638
rect 491062 149636 491083 149640
rect 495802 149638 495894 149698
rect 495888 149636 495894 149638
rect 495958 149636 495964 149700
rect 503504 149698 503510 149700
rect 503438 149638 503510 149698
rect 503574 149696 503595 149700
rect 503590 149640 503595 149696
rect 503504 149636 503510 149638
rect 503574 149636 503595 149640
rect 488257 149635 488323 149636
rect 491017 149635 491083 149636
rect 495893 149635 495959 149636
rect 503529 149635 503595 149636
rect 48313 149564 48379 149565
rect 50797 149564 50863 149565
rect 56041 149564 56107 149565
rect 58525 149564 58591 149565
rect 48288 149562 48294 149564
rect 48222 149502 48294 149562
rect 48358 149560 48379 149564
rect 50736 149562 50742 149564
rect 48374 149504 48379 149560
rect 48288 149500 48294 149502
rect 48358 149500 48379 149504
rect 50706 149502 50742 149562
rect 50806 149560 50863 149564
rect 50858 149504 50863 149560
rect 50736 149500 50742 149502
rect 50806 149500 50863 149504
rect 56040 149500 56046 149564
rect 56110 149562 56116 149564
rect 58488 149562 58494 149564
rect 56110 149502 56198 149562
rect 58434 149502 58494 149562
rect 58558 149560 58591 149564
rect 58586 149504 58591 149560
rect 56110 149500 56116 149502
rect 58488 149500 58494 149502
rect 58558 149500 58591 149504
rect 48313 149499 48379 149500
rect 50797 149499 50863 149500
rect 56041 149499 56107 149500
rect 58525 149499 58591 149500
rect 60641 149564 60707 149565
rect 60641 149560 60670 149564
rect 60734 149562 60740 149564
rect 60641 149504 60646 149560
rect 60641 149500 60670 149504
rect 60734 149502 60798 149562
rect 60734 149500 60740 149502
rect 71000 149500 71006 149564
rect 71070 149562 71076 149564
rect 71221 149562 71287 149565
rect 73613 149564 73679 149565
rect 83549 149564 83615 149565
rect 93485 149564 93551 149565
rect 98545 149564 98611 149565
rect 103513 149564 103579 149565
rect 113449 149564 113515 149565
rect 73584 149562 73590 149564
rect 71070 149560 71287 149562
rect 71070 149504 71226 149560
rect 71282 149504 71287 149560
rect 71070 149502 71287 149504
rect 73522 149502 73590 149562
rect 73654 149560 73679 149564
rect 83512 149562 83518 149564
rect 73674 149504 73679 149560
rect 71070 149500 71076 149502
rect 60641 149499 60707 149500
rect 71221 149499 71287 149502
rect 73584 149500 73590 149502
rect 73654 149500 73679 149504
rect 83458 149502 83518 149562
rect 83582 149560 83615 149564
rect 93440 149562 93446 149564
rect 83610 149504 83615 149560
rect 83512 149500 83518 149502
rect 83582 149500 83615 149504
rect 93394 149502 93446 149562
rect 93510 149560 93551 149564
rect 98472 149562 98478 149564
rect 93546 149504 93551 149560
rect 93440 149500 93446 149502
rect 93510 149500 93551 149504
rect 98454 149502 98478 149562
rect 98472 149500 98478 149502
rect 98542 149560 98611 149564
rect 103504 149562 103510 149564
rect 98542 149504 98550 149560
rect 98606 149504 98611 149560
rect 98542 149500 98611 149504
rect 103422 149502 103510 149562
rect 103504 149500 103510 149502
rect 103574 149500 103580 149564
rect 113432 149562 113438 149564
rect 113358 149502 113438 149562
rect 113502 149560 113515 149564
rect 113510 149504 113515 149560
rect 113432 149500 113438 149502
rect 113502 149500 113515 149504
rect 73613 149499 73679 149500
rect 83549 149499 83615 149500
rect 93485 149499 93551 149500
rect 98545 149499 98611 149500
rect 103513 149499 103579 149500
rect 113449 149499 113515 149500
rect 115841 149564 115907 149565
rect 120901 149564 120967 149565
rect 115841 149560 115886 149564
rect 115950 149562 115956 149564
rect 115841 149504 115846 149560
rect 115841 149500 115886 149504
rect 115950 149502 115998 149562
rect 120901 149560 120918 149564
rect 120982 149562 120988 149564
rect 438209 149562 438275 149565
rect 441760 149562 441766 149564
rect 120901 149504 120906 149560
rect 115950 149500 115956 149502
rect 120901 149500 120918 149504
rect 120982 149502 121058 149562
rect 438209 149560 441766 149562
rect 438209 149504 438214 149560
rect 438270 149504 441766 149560
rect 438209 149502 441766 149504
rect 120982 149500 120988 149502
rect 115841 149499 115907 149500
rect 120901 149499 120967 149500
rect 438209 149499 438275 149502
rect 441760 149500 441766 149502
rect 441830 149500 441836 149564
rect 455904 149500 455910 149564
rect 455974 149562 455980 149564
rect 456793 149562 456859 149565
rect 463509 149564 463575 149565
rect 465993 149564 466059 149565
rect 468293 149564 468359 149565
rect 455974 149560 456859 149562
rect 455974 149504 456798 149560
rect 456854 149504 456859 149560
rect 455974 149502 456859 149504
rect 455974 149500 455980 149502
rect 456793 149499 456859 149502
rect 461072 149500 461078 149564
rect 461142 149500 461148 149564
rect 463509 149560 463526 149564
rect 463590 149562 463596 149564
rect 465968 149562 465974 149564
rect 463509 149504 463514 149560
rect 463509 149500 463526 149504
rect 463590 149502 463666 149562
rect 465902 149502 465974 149562
rect 466038 149560 466059 149564
rect 468280 149562 468286 149564
rect 466054 149504 466059 149560
rect 463590 149500 463596 149502
rect 465968 149500 465974 149502
rect 466038 149500 466059 149504
rect 468202 149502 468286 149562
rect 468350 149560 468359 149564
rect 468354 149504 468359 149560
rect 468280 149500 468286 149502
rect 468350 149500 468359 149504
rect 406837 149290 406903 149293
rect 461080 149290 461140 149500
rect 463509 149499 463575 149500
rect 465993 149499 466059 149500
rect 468293 149499 468359 149500
rect 470961 149564 471027 149565
rect 505921 149564 505987 149565
rect 508497 149564 508563 149565
rect 510981 149564 511047 149565
rect 515857 149564 515923 149565
rect 518433 149564 518499 149565
rect 470961 149560 471006 149564
rect 471070 149562 471076 149564
rect 470961 149504 470966 149560
rect 470961 149500 471006 149504
rect 471070 149502 471118 149562
rect 505921 149560 505958 149564
rect 506022 149562 506028 149564
rect 505921 149504 505926 149560
rect 471070 149500 471076 149502
rect 505921 149500 505958 149504
rect 506022 149502 506078 149562
rect 508497 149560 508542 149564
rect 508606 149562 508612 149564
rect 508497 149504 508502 149560
rect 506022 149500 506028 149502
rect 508497 149500 508542 149504
rect 508606 149502 508654 149562
rect 510981 149560 510990 149564
rect 511054 149562 511060 149564
rect 510981 149504 510986 149560
rect 508606 149500 508612 149502
rect 510981 149500 510990 149504
rect 511054 149502 511138 149562
rect 515857 149560 515886 149564
rect 515950 149562 515956 149564
rect 515857 149504 515862 149560
rect 511054 149500 511060 149502
rect 515857 149500 515886 149504
rect 515950 149502 516014 149562
rect 518433 149560 518470 149564
rect 518534 149562 518540 149564
rect 518433 149504 518438 149560
rect 515950 149500 515956 149502
rect 518433 149500 518470 149504
rect 518534 149502 518590 149562
rect 518534 149500 518540 149502
rect 470961 149499 471027 149500
rect 505921 149499 505987 149500
rect 508497 149499 508563 149500
rect 510981 149499 511047 149500
rect 515857 149499 515923 149500
rect 518433 149499 518499 149500
rect 406837 149288 461140 149290
rect 406837 149232 406842 149288
rect 406898 149232 461140 149288
rect 406837 149230 461140 149232
rect 406837 149227 406903 149230
rect 414933 149154 414999 149157
rect 476062 149154 476068 149156
rect 414933 149152 476068 149154
rect 414933 149096 414938 149152
rect 414994 149096 476068 149152
rect 414933 149094 476068 149096
rect 414933 149091 414999 149094
rect 476062 149092 476068 149094
rect 476132 149092 476138 149156
rect 53649 149020 53715 149021
rect 76097 149020 76163 149021
rect 86033 149020 86099 149021
rect 53598 149018 53604 149020
rect 53558 148958 53604 149018
rect 53668 149016 53715 149020
rect 76046 149018 76052 149020
rect 53710 148960 53715 149016
rect 53598 148956 53604 148958
rect 53668 148956 53715 148960
rect 76006 148958 76052 149018
rect 76116 149016 76163 149020
rect 85982 149018 85988 149020
rect 76158 148960 76163 149016
rect 76046 148956 76052 148958
rect 76116 148956 76163 148960
rect 85942 148958 85988 149018
rect 86052 149016 86099 149020
rect 86094 148960 86099 149016
rect 85982 148956 85988 148958
rect 86052 148956 86099 148960
rect 123334 148956 123340 149020
rect 123404 149018 123410 149020
rect 183185 149018 183251 149021
rect 123404 149016 183251 149018
rect 123404 148960 183190 149016
rect 183246 148960 183251 149016
rect 123404 148958 183251 148960
rect 123404 148956 123410 148958
rect 53649 148955 53715 148956
rect 76097 148955 76163 148956
rect 86033 148955 86099 148956
rect 183185 148955 183251 148958
rect 513373 149020 513439 149021
rect 520917 149020 520983 149021
rect 523309 149020 523375 149021
rect 525885 149020 525951 149021
rect 513373 149016 513420 149020
rect 513484 149018 513490 149020
rect 513373 148960 513378 149016
rect 513373 148956 513420 148960
rect 513484 148958 513530 149018
rect 520917 149016 520964 149020
rect 521028 149018 521034 149020
rect 520917 148960 520922 149016
rect 513484 148956 513490 148958
rect 520917 148956 520964 148960
rect 521028 148958 521074 149018
rect 523309 149016 523356 149020
rect 523420 149018 523426 149020
rect 523309 148960 523314 149016
rect 521028 148956 521034 148958
rect 523309 148956 523356 148960
rect 523420 148958 523466 149018
rect 525885 149016 525932 149020
rect 525996 149018 526002 149020
rect 525885 148960 525890 149016
rect 523420 148956 523426 148958
rect 525885 148956 525932 148960
rect 525996 148958 526042 149018
rect 525996 148956 526002 148958
rect 513373 148955 513439 148956
rect 520917 148955 520983 148956
rect 523309 148955 523375 148956
rect 525885 148955 525951 148956
rect 125910 148820 125916 148884
rect 125980 148882 125986 148884
rect 183369 148882 183435 148885
rect 125980 148880 183435 148882
rect 125980 148824 183374 148880
rect 183430 148824 183435 148880
rect 125980 148822 183435 148824
rect 125980 148820 125986 148822
rect 183369 148819 183435 148822
rect 459461 148748 459527 148749
rect 459461 148746 459508 148748
rect 459416 148744 459508 148746
rect 459416 148688 459466 148744
rect 459416 148686 459508 148688
rect 459461 148684 459508 148686
rect 459572 148684 459578 148748
rect 459461 148683 459527 148684
rect 419942 148276 419948 148340
rect 420012 148338 420018 148340
rect 459461 148338 459527 148341
rect 420012 148336 459527 148338
rect 420012 148280 459466 148336
rect 459522 148280 459527 148336
rect 420012 148278 459527 148280
rect 420012 148276 420018 148278
rect 459461 148275 459527 148278
rect 35893 147660 35959 147661
rect 36997 147660 37063 147661
rect 38101 147660 38167 147661
rect 39573 147660 39639 147661
rect 43069 147660 43135 147661
rect 44173 147660 44239 147661
rect 45277 147660 45343 147661
rect 46565 147660 46631 147661
rect 47669 147660 47735 147661
rect 48681 147660 48747 147661
rect 50153 147660 50219 147661
rect 51441 147660 51507 147661
rect 35893 147656 35940 147660
rect 36004 147658 36010 147660
rect 35893 147600 35898 147656
rect 35893 147596 35940 147600
rect 36004 147598 36050 147658
rect 36997 147656 37044 147660
rect 37108 147658 37114 147660
rect 36997 147600 37002 147656
rect 36004 147596 36010 147598
rect 36997 147596 37044 147600
rect 37108 147598 37154 147658
rect 38101 147656 38148 147660
rect 38212 147658 38218 147660
rect 38101 147600 38106 147656
rect 37108 147596 37114 147598
rect 38101 147596 38148 147600
rect 38212 147598 38258 147658
rect 39573 147656 39620 147660
rect 39684 147658 39690 147660
rect 39573 147600 39578 147656
rect 38212 147596 38218 147598
rect 39573 147596 39620 147600
rect 39684 147598 39730 147658
rect 43069 147656 43116 147660
rect 43180 147658 43186 147660
rect 43069 147600 43074 147656
rect 39684 147596 39690 147598
rect 43069 147596 43116 147600
rect 43180 147598 43226 147658
rect 44173 147656 44220 147660
rect 44284 147658 44290 147660
rect 44173 147600 44178 147656
rect 43180 147596 43186 147598
rect 44173 147596 44220 147600
rect 44284 147598 44330 147658
rect 45277 147656 45324 147660
rect 45388 147658 45394 147660
rect 45277 147600 45282 147656
rect 44284 147596 44290 147598
rect 45277 147596 45324 147600
rect 45388 147598 45434 147658
rect 46565 147656 46612 147660
rect 46676 147658 46682 147660
rect 46565 147600 46570 147656
rect 45388 147596 45394 147598
rect 46565 147596 46612 147600
rect 46676 147598 46722 147658
rect 47669 147656 47716 147660
rect 47780 147658 47786 147660
rect 48630 147658 48636 147660
rect 47669 147600 47674 147656
rect 46676 147596 46682 147598
rect 47669 147596 47716 147600
rect 47780 147598 47826 147658
rect 48590 147598 48636 147658
rect 48700 147656 48747 147660
rect 50102 147658 50108 147660
rect 48742 147600 48747 147656
rect 47780 147596 47786 147598
rect 48630 147596 48636 147598
rect 48700 147596 48747 147600
rect 50062 147598 50108 147658
rect 50172 147656 50219 147660
rect 51390 147658 51396 147660
rect 50214 147600 50219 147656
rect 50102 147596 50108 147598
rect 50172 147596 50219 147600
rect 51350 147598 51396 147658
rect 51460 147656 51507 147660
rect 51502 147600 51507 147656
rect 51390 147596 51396 147598
rect 51460 147596 51507 147600
rect 35893 147595 35959 147596
rect 36997 147595 37063 147596
rect 38101 147595 38167 147596
rect 39573 147595 39639 147596
rect 43069 147595 43135 147596
rect 44173 147595 44239 147596
rect 45277 147595 45343 147596
rect 46565 147595 46631 147596
rect 47669 147595 47735 147596
rect 48681 147595 48747 147596
rect 50153 147595 50219 147596
rect 51441 147595 51507 147596
rect 52269 147660 52335 147661
rect 53373 147660 53439 147661
rect 52269 147656 52316 147660
rect 52380 147658 52386 147660
rect 52269 147600 52274 147656
rect 52269 147596 52316 147600
rect 52380 147598 52426 147658
rect 53373 147656 53420 147660
rect 53484 147658 53490 147660
rect 54017 147658 54083 147661
rect 56041 147660 56107 147661
rect 58065 147660 58131 147661
rect 59537 147660 59603 147661
rect 54518 147658 54524 147660
rect 53373 147600 53378 147656
rect 52380 147596 52386 147598
rect 53373 147596 53420 147600
rect 53484 147598 53530 147658
rect 54017 147656 54524 147658
rect 54017 147600 54022 147656
rect 54078 147600 54524 147656
rect 54017 147598 54524 147600
rect 53484 147596 53490 147598
rect 52269 147595 52335 147596
rect 53373 147595 53439 147596
rect 54017 147595 54083 147598
rect 54518 147596 54524 147598
rect 54588 147596 54594 147660
rect 55990 147658 55996 147660
rect 55950 147598 55996 147658
rect 56060 147656 56107 147660
rect 58014 147658 58020 147660
rect 56102 147600 56107 147656
rect 55990 147596 55996 147598
rect 56060 147596 56107 147600
rect 57974 147598 58020 147658
rect 58084 147656 58131 147660
rect 59486 147658 59492 147660
rect 58126 147600 58131 147656
rect 58014 147596 58020 147598
rect 58084 147596 58131 147600
rect 59446 147598 59492 147658
rect 59556 147656 59603 147660
rect 59598 147600 59603 147656
rect 59486 147596 59492 147598
rect 59556 147596 59603 147600
rect 56041 147595 56107 147596
rect 58065 147595 58131 147596
rect 59537 147595 59603 147596
rect 61653 147660 61719 147661
rect 62757 147660 62823 147661
rect 63585 147660 63651 147661
rect 61653 147656 61700 147660
rect 61764 147658 61770 147660
rect 61653 147600 61658 147656
rect 61653 147596 61700 147600
rect 61764 147598 61810 147658
rect 62757 147656 62804 147660
rect 62868 147658 62874 147660
rect 63534 147658 63540 147660
rect 62757 147600 62762 147656
rect 61764 147596 61770 147598
rect 62757 147596 62804 147600
rect 62868 147598 62914 147658
rect 63494 147598 63540 147658
rect 63604 147656 63651 147660
rect 63646 147600 63651 147656
rect 62868 147596 62874 147598
rect 63534 147596 63540 147598
rect 63604 147596 63651 147600
rect 61653 147595 61719 147596
rect 62757 147595 62823 147596
rect 63585 147595 63651 147596
rect 63861 147660 63927 147661
rect 65149 147660 65215 147661
rect 66161 147660 66227 147661
rect 66345 147660 66411 147661
rect 67633 147660 67699 147661
rect 63861 147656 63908 147660
rect 63972 147658 63978 147660
rect 63861 147600 63866 147656
rect 63861 147596 63908 147600
rect 63972 147598 64018 147658
rect 65149 147656 65196 147660
rect 65260 147658 65266 147660
rect 66110 147658 66116 147660
rect 65149 147600 65154 147656
rect 63972 147596 63978 147598
rect 65149 147596 65196 147600
rect 65260 147598 65306 147658
rect 66070 147598 66116 147658
rect 66180 147656 66227 147660
rect 66222 147600 66227 147656
rect 65260 147596 65266 147598
rect 66110 147596 66116 147598
rect 66180 147596 66227 147600
rect 66294 147596 66300 147660
rect 66364 147658 66411 147660
rect 67582 147658 67588 147660
rect 66364 147656 66456 147658
rect 66406 147600 66456 147656
rect 66364 147598 66456 147600
rect 67542 147598 67588 147658
rect 67652 147656 67699 147660
rect 67694 147600 67699 147656
rect 66364 147596 66411 147598
rect 67582 147596 67588 147598
rect 67652 147596 67699 147600
rect 68134 147596 68140 147660
rect 68204 147658 68210 147660
rect 68277 147658 68343 147661
rect 68204 147656 68343 147658
rect 68204 147600 68282 147656
rect 68338 147600 68343 147656
rect 68204 147598 68343 147600
rect 68204 147596 68210 147598
rect 63861 147595 63927 147596
rect 65149 147595 65215 147596
rect 66161 147595 66227 147596
rect 66345 147595 66411 147596
rect 67633 147595 67699 147596
rect 68277 147595 68343 147598
rect 68461 147658 68527 147661
rect 69749 147660 69815 147661
rect 72141 147660 72207 147661
rect 73245 147660 73311 147661
rect 68686 147658 68692 147660
rect 68461 147656 68692 147658
rect 68461 147600 68466 147656
rect 68522 147600 68692 147656
rect 68461 147598 68692 147600
rect 68461 147595 68527 147598
rect 68686 147596 68692 147598
rect 68756 147596 68762 147660
rect 69749 147656 69796 147660
rect 69860 147658 69866 147660
rect 69749 147600 69754 147656
rect 69749 147596 69796 147600
rect 69860 147598 69906 147658
rect 72141 147656 72188 147660
rect 72252 147658 72258 147660
rect 72141 147600 72146 147656
rect 69860 147596 69866 147598
rect 72141 147596 72188 147600
rect 72252 147598 72298 147658
rect 73245 147656 73292 147660
rect 73356 147658 73362 147660
rect 73705 147658 73771 147661
rect 75637 147660 75703 147661
rect 76925 147660 76991 147661
rect 78029 147660 78095 147661
rect 78489 147660 78555 147661
rect 74390 147658 74396 147660
rect 73245 147600 73250 147656
rect 72252 147596 72258 147598
rect 73245 147596 73292 147600
rect 73356 147598 73402 147658
rect 73705 147656 74396 147658
rect 73705 147600 73710 147656
rect 73766 147600 74396 147656
rect 73705 147598 74396 147600
rect 73356 147596 73362 147598
rect 69749 147595 69815 147596
rect 72141 147595 72207 147596
rect 73245 147595 73311 147596
rect 73705 147595 73771 147598
rect 74390 147596 74396 147598
rect 74460 147596 74466 147660
rect 75637 147656 75684 147660
rect 75748 147658 75754 147660
rect 75637 147600 75642 147656
rect 75637 147596 75684 147600
rect 75748 147598 75794 147658
rect 76925 147656 76972 147660
rect 77036 147658 77042 147660
rect 76925 147600 76930 147656
rect 75748 147596 75754 147598
rect 76925 147596 76972 147600
rect 77036 147598 77082 147658
rect 78029 147656 78076 147660
rect 78140 147658 78146 147660
rect 78438 147658 78444 147660
rect 78029 147600 78034 147656
rect 77036 147596 77042 147598
rect 78029 147596 78076 147600
rect 78140 147598 78186 147658
rect 78398 147598 78444 147658
rect 78508 147656 78555 147660
rect 78550 147600 78555 147656
rect 78140 147596 78146 147598
rect 78438 147596 78444 147598
rect 78508 147596 78555 147600
rect 75637 147595 75703 147596
rect 76925 147595 76991 147596
rect 78029 147595 78095 147596
rect 78489 147595 78555 147596
rect 79133 147660 79199 147661
rect 81065 147660 81131 147661
rect 88241 147660 88307 147661
rect 91001 147660 91067 147661
rect 95969 147660 96035 147661
rect 100937 147660 101003 147661
rect 106089 147660 106155 147661
rect 79133 147656 79180 147660
rect 79244 147658 79250 147660
rect 81014 147658 81020 147660
rect 79133 147600 79138 147656
rect 79133 147596 79180 147600
rect 79244 147598 79290 147658
rect 80974 147598 81020 147658
rect 81084 147656 81131 147660
rect 88190 147658 88196 147660
rect 81126 147600 81131 147656
rect 79244 147596 79250 147598
rect 81014 147596 81020 147598
rect 81084 147596 81131 147600
rect 88150 147598 88196 147658
rect 88260 147656 88307 147660
rect 90950 147658 90956 147660
rect 88302 147600 88307 147656
rect 88190 147596 88196 147598
rect 88260 147596 88307 147600
rect 90910 147598 90956 147658
rect 91020 147656 91067 147660
rect 95918 147658 95924 147660
rect 91062 147600 91067 147656
rect 90950 147596 90956 147598
rect 91020 147596 91067 147600
rect 95878 147598 95924 147658
rect 95988 147656 96035 147660
rect 100886 147658 100892 147660
rect 96030 147600 96035 147656
rect 95918 147596 95924 147598
rect 95988 147596 96035 147600
rect 100846 147598 100892 147658
rect 100956 147656 101003 147660
rect 106038 147658 106044 147660
rect 100998 147600 101003 147656
rect 100886 147596 100892 147598
rect 100956 147596 101003 147600
rect 105998 147598 106044 147658
rect 106108 147656 106155 147660
rect 106150 147600 106155 147656
rect 106038 147596 106044 147598
rect 106108 147596 106155 147600
rect 108614 147596 108620 147660
rect 108684 147658 108690 147660
rect 108849 147658 108915 147661
rect 108684 147656 108915 147658
rect 108684 147600 108854 147656
rect 108910 147600 108915 147656
rect 108684 147598 108915 147600
rect 108684 147596 108690 147598
rect 79133 147595 79199 147596
rect 81065 147595 81131 147596
rect 88241 147595 88307 147596
rect 91001 147595 91067 147596
rect 95969 147595 96035 147596
rect 100937 147595 101003 147596
rect 106089 147595 106155 147596
rect 108849 147595 108915 147598
rect 111006 147596 111012 147660
rect 111076 147658 111082 147660
rect 111609 147658 111675 147661
rect 111076 147656 111675 147658
rect 111076 147600 111614 147656
rect 111670 147600 111675 147656
rect 111076 147598 111675 147600
rect 111076 147596 111082 147598
rect 111609 147595 111675 147598
rect 436093 147660 436159 147661
rect 437013 147660 437079 147661
rect 437933 147660 437999 147661
rect 439589 147660 439655 147661
rect 443085 147660 443151 147661
rect 444189 147660 444255 147661
rect 445293 147660 445359 147661
rect 446397 147660 446463 147661
rect 436093 147656 436140 147660
rect 436204 147658 436210 147660
rect 436093 147600 436098 147656
rect 436093 147596 436140 147600
rect 436204 147598 436250 147658
rect 437013 147656 437060 147660
rect 437124 147658 437130 147660
rect 437013 147600 437018 147656
rect 436204 147596 436210 147598
rect 437013 147596 437060 147600
rect 437124 147598 437170 147658
rect 437933 147656 437980 147660
rect 438044 147658 438050 147660
rect 437933 147600 437938 147656
rect 437124 147596 437130 147598
rect 437933 147596 437980 147600
rect 438044 147598 438090 147658
rect 439589 147656 439636 147660
rect 439700 147658 439706 147660
rect 439589 147600 439594 147656
rect 438044 147596 438050 147598
rect 439589 147596 439636 147600
rect 439700 147598 439746 147658
rect 443085 147656 443132 147660
rect 443196 147658 443202 147660
rect 443085 147600 443090 147656
rect 439700 147596 439706 147598
rect 443085 147596 443132 147600
rect 443196 147598 443242 147658
rect 444189 147656 444236 147660
rect 444300 147658 444306 147660
rect 444189 147600 444194 147656
rect 443196 147596 443202 147598
rect 444189 147596 444236 147600
rect 444300 147598 444346 147658
rect 445293 147656 445340 147660
rect 445404 147658 445410 147660
rect 445293 147600 445298 147656
rect 444300 147596 444306 147598
rect 445293 147596 445340 147600
rect 445404 147598 445450 147658
rect 446397 147656 446444 147660
rect 446508 147658 446514 147660
rect 447133 147658 447199 147661
rect 448237 147660 448303 147661
rect 447358 147658 447364 147660
rect 446397 147600 446402 147656
rect 445404 147596 445410 147598
rect 446397 147596 446444 147600
rect 446508 147598 446554 147658
rect 447133 147656 447364 147658
rect 447133 147600 447138 147656
rect 447194 147600 447364 147656
rect 447133 147598 447364 147600
rect 446508 147596 446514 147598
rect 436093 147595 436159 147596
rect 437013 147595 437079 147596
rect 437933 147595 437999 147596
rect 439589 147595 439655 147596
rect 443085 147595 443151 147596
rect 444189 147595 444255 147596
rect 445293 147595 445359 147596
rect 446397 147595 446463 147596
rect 447133 147595 447199 147598
rect 447358 147596 447364 147598
rect 447428 147596 447434 147660
rect 448237 147656 448284 147660
rect 448348 147658 448354 147660
rect 448513 147658 448579 147661
rect 448646 147658 448652 147660
rect 448237 147600 448242 147656
rect 448237 147596 448284 147600
rect 448348 147598 448394 147658
rect 448513 147656 448652 147658
rect 448513 147600 448518 147656
rect 448574 147600 448652 147656
rect 448513 147598 448652 147600
rect 448348 147596 448354 147598
rect 448237 147595 448303 147596
rect 448513 147595 448579 147598
rect 448646 147596 448652 147598
rect 448716 147596 448722 147660
rect 449893 147658 449959 147661
rect 450629 147660 450695 147661
rect 451273 147660 451339 147661
rect 450118 147658 450124 147660
rect 449893 147656 450124 147658
rect 449893 147600 449898 147656
rect 449954 147600 450124 147656
rect 449893 147598 450124 147600
rect 449893 147595 449959 147598
rect 450118 147596 450124 147598
rect 450188 147596 450194 147660
rect 450629 147656 450676 147660
rect 450740 147658 450746 147660
rect 450629 147600 450634 147656
rect 450629 147596 450676 147600
rect 450740 147598 450786 147658
rect 450740 147596 450746 147598
rect 451222 147596 451228 147660
rect 451292 147658 451339 147660
rect 451292 147656 451384 147658
rect 451334 147600 451384 147656
rect 451292 147598 451384 147600
rect 451292 147596 451339 147598
rect 452326 147596 452332 147660
rect 452396 147658 452402 147660
rect 452561 147658 452627 147661
rect 453389 147660 453455 147661
rect 453573 147660 453639 147661
rect 454585 147660 454651 147661
rect 453389 147658 453436 147660
rect 452396 147656 452627 147658
rect 452396 147600 452566 147656
rect 452622 147600 452627 147656
rect 452396 147598 452627 147600
rect 453344 147656 453436 147658
rect 453344 147600 453394 147656
rect 453344 147598 453436 147600
rect 452396 147596 452402 147598
rect 450629 147595 450695 147596
rect 451273 147595 451339 147596
rect 452561 147595 452627 147598
rect 453389 147596 453436 147598
rect 453500 147596 453506 147660
rect 453573 147656 453620 147660
rect 453684 147658 453690 147660
rect 454534 147658 454540 147660
rect 453573 147600 453578 147656
rect 453573 147596 453620 147600
rect 453684 147598 453730 147658
rect 454494 147598 454540 147658
rect 454604 147656 454651 147660
rect 454646 147600 454651 147656
rect 453684 147596 453690 147598
rect 454534 147596 454540 147598
rect 454604 147596 454651 147600
rect 453389 147595 453455 147596
rect 453573 147595 453639 147596
rect 454585 147595 454651 147596
rect 455965 147660 456031 147661
rect 458357 147660 458423 147661
rect 461669 147660 461735 147661
rect 462773 147660 462839 147661
rect 463877 147660 463943 147661
rect 465165 147660 465231 147661
rect 466269 147660 466335 147661
rect 467557 147660 467623 147661
rect 468661 147660 468727 147661
rect 469765 147660 469831 147661
rect 471053 147660 471119 147661
rect 472157 147660 472223 147661
rect 473353 147660 473419 147661
rect 455965 147656 456012 147660
rect 456076 147658 456082 147660
rect 455965 147600 455970 147656
rect 455965 147596 456012 147600
rect 456076 147598 456122 147658
rect 458357 147656 458404 147660
rect 458468 147658 458474 147660
rect 458357 147600 458362 147656
rect 456076 147596 456082 147598
rect 458357 147596 458404 147600
rect 458468 147598 458514 147658
rect 461669 147656 461716 147660
rect 461780 147658 461786 147660
rect 461669 147600 461674 147656
rect 458468 147596 458474 147598
rect 461669 147596 461716 147600
rect 461780 147598 461826 147658
rect 462773 147656 462820 147660
rect 462884 147658 462890 147660
rect 462773 147600 462778 147656
rect 461780 147596 461786 147598
rect 462773 147596 462820 147600
rect 462884 147598 462930 147658
rect 463877 147656 463924 147660
rect 463988 147658 463994 147660
rect 463877 147600 463882 147656
rect 462884 147596 462890 147598
rect 463877 147596 463924 147600
rect 463988 147598 464034 147658
rect 465165 147656 465212 147660
rect 465276 147658 465282 147660
rect 465165 147600 465170 147656
rect 463988 147596 463994 147598
rect 465165 147596 465212 147600
rect 465276 147598 465322 147658
rect 466269 147656 466316 147660
rect 466380 147658 466386 147660
rect 466269 147600 466274 147656
rect 465276 147596 465282 147598
rect 466269 147596 466316 147600
rect 466380 147598 466426 147658
rect 467557 147656 467604 147660
rect 467668 147658 467674 147660
rect 467557 147600 467562 147656
rect 466380 147596 466386 147598
rect 467557 147596 467604 147600
rect 467668 147598 467714 147658
rect 468661 147656 468708 147660
rect 468772 147658 468778 147660
rect 468661 147600 468666 147656
rect 467668 147596 467674 147598
rect 468661 147596 468708 147600
rect 468772 147598 468818 147658
rect 469765 147656 469812 147660
rect 469876 147658 469882 147660
rect 469765 147600 469770 147656
rect 468772 147596 468778 147598
rect 469765 147596 469812 147600
rect 469876 147598 469922 147658
rect 471053 147656 471100 147660
rect 471164 147658 471170 147660
rect 471053 147600 471058 147656
rect 469876 147596 469882 147598
rect 471053 147596 471100 147600
rect 471164 147598 471210 147658
rect 472157 147656 472204 147660
rect 472268 147658 472274 147660
rect 473302 147658 473308 147660
rect 472157 147600 472162 147656
rect 471164 147596 471170 147598
rect 472157 147596 472204 147600
rect 472268 147598 472314 147658
rect 473262 147598 473308 147658
rect 473372 147656 473419 147660
rect 473414 147600 473419 147656
rect 472268 147596 472274 147598
rect 473302 147596 473308 147598
rect 473372 147596 473419 147600
rect 455965 147595 456031 147596
rect 458357 147595 458423 147596
rect 461669 147595 461735 147596
rect 462773 147595 462839 147596
rect 463877 147595 463943 147596
rect 465165 147595 465231 147596
rect 466269 147595 466335 147596
rect 467557 147595 467623 147596
rect 468661 147595 468727 147596
rect 469765 147595 469831 147596
rect 471053 147595 471119 147596
rect 472157 147595 472223 147596
rect 473353 147595 473419 147596
rect 474089 147658 474155 147661
rect 476941 147660 477007 147661
rect 478045 147660 478111 147661
rect 474406 147658 474412 147660
rect 474089 147656 474412 147658
rect 474089 147600 474094 147656
rect 474150 147600 474412 147656
rect 474089 147598 474412 147600
rect 474089 147595 474155 147598
rect 474406 147596 474412 147598
rect 474476 147596 474482 147660
rect 476941 147656 476988 147660
rect 477052 147658 477058 147660
rect 476941 147600 476946 147656
rect 476941 147596 476988 147600
rect 477052 147598 477098 147658
rect 478045 147656 478092 147660
rect 478156 147658 478162 147660
rect 478045 147600 478050 147656
rect 477052 147596 477058 147598
rect 478045 147596 478092 147600
rect 478156 147598 478202 147658
rect 478156 147596 478162 147598
rect 476941 147595 477007 147596
rect 478045 147595 478111 147596
rect 18638 147460 18644 147524
rect 18708 147522 18714 147524
rect 41822 147522 41828 147524
rect 18708 147462 41828 147522
rect 18708 147460 18714 147462
rect 41822 147460 41828 147462
rect 41892 147460 41898 147524
rect 60641 147522 60707 147525
rect 75821 147522 75887 147525
rect 60641 147520 75887 147522
rect 60641 147464 60646 147520
rect 60702 147464 75826 147520
rect 75882 147464 75887 147520
rect 60641 147462 75887 147464
rect 60641 147459 60707 147462
rect 75821 147459 75887 147462
rect 118550 147460 118556 147524
rect 118620 147522 118626 147524
rect 156781 147522 156847 147525
rect 118620 147520 156847 147522
rect 118620 147464 156786 147520
rect 156842 147464 156847 147520
rect 118620 147462 156847 147464
rect 118620 147460 118626 147462
rect 156781 147459 156847 147462
rect 392577 147522 392643 147525
rect 500902 147522 500908 147524
rect 392577 147520 500908 147522
rect 392577 147464 392582 147520
rect 392638 147464 500908 147520
rect 392577 147462 500908 147464
rect 392577 147459 392643 147462
rect 500902 147460 500908 147462
rect 500972 147460 500978 147524
rect 19425 147386 19491 147389
rect 40534 147386 40540 147388
rect 19425 147384 40540 147386
rect 19425 147328 19430 147384
rect 19486 147328 40540 147384
rect 19425 147326 40540 147328
rect 19425 147323 19491 147326
rect 40534 147324 40540 147326
rect 40604 147324 40610 147388
rect 61142 147324 61148 147388
rect 61212 147386 61218 147388
rect 180149 147386 180215 147389
rect 61212 147384 180215 147386
rect 61212 147328 180154 147384
rect 180210 147328 180215 147384
rect 61212 147326 180215 147328
rect 61212 147324 61218 147326
rect 180149 147323 180215 147326
rect 388437 147386 388503 147389
rect 493358 147386 493364 147388
rect 388437 147384 493364 147386
rect 388437 147328 388442 147384
rect 388498 147328 493364 147384
rect 388437 147326 493364 147328
rect 388437 147323 388503 147326
rect 493358 147324 493364 147326
rect 493428 147324 493434 147388
rect 19517 147250 19583 147253
rect 56910 147250 56916 147252
rect 19517 147248 56916 147250
rect 19517 147192 19522 147248
rect 19578 147192 56916 147248
rect 19517 147190 56916 147192
rect 19517 147187 19583 147190
rect 56910 147188 56916 147190
rect 56980 147250 56986 147252
rect 70393 147250 70459 147253
rect 56980 147248 70459 147250
rect 56980 147192 70398 147248
rect 70454 147192 70459 147248
rect 56980 147190 70459 147192
rect 56980 147188 56986 147190
rect 70393 147187 70459 147190
rect 71037 147252 71103 147253
rect 71037 147248 71084 147252
rect 71148 147250 71154 147252
rect 71037 147192 71042 147248
rect 71037 147188 71084 147192
rect 71148 147190 71194 147250
rect 71148 147188 71154 147190
rect 419390 147188 419396 147252
rect 419460 147250 419466 147252
rect 440049 147250 440115 147253
rect 419460 147248 440115 147250
rect 419460 147192 440054 147248
rect 440110 147192 440115 147248
rect 419460 147190 440115 147192
rect 419460 147188 419466 147190
rect 71037 147187 71103 147188
rect 440049 147187 440115 147190
rect 440233 147250 440299 147253
rect 473486 147250 473492 147252
rect 440233 147248 473492 147250
rect 440233 147192 440238 147248
rect 440294 147192 473492 147248
rect 440233 147190 473492 147192
rect 440233 147187 440299 147190
rect 473486 147188 473492 147190
rect 473556 147188 473562 147252
rect 418061 147114 418127 147117
rect 418705 147114 418771 147117
rect 456926 147114 456932 147116
rect 418061 147112 456932 147114
rect 418061 147056 418066 147112
rect 418122 147056 418710 147112
rect 418766 147056 456932 147112
rect 418061 147054 456932 147056
rect 418061 147051 418127 147054
rect 418705 147051 418771 147054
rect 456926 147052 456932 147054
rect 456996 147052 457002 147116
rect 479190 147114 479196 147116
rect 460890 147054 479196 147114
rect 417785 146978 417851 146981
rect 418797 146978 418863 146981
rect 460606 146978 460612 146980
rect 417785 146976 460612 146978
rect 417785 146920 417790 146976
rect 417846 146920 418802 146976
rect 418858 146920 460612 146976
rect 417785 146918 460612 146920
rect 417785 146915 417851 146918
rect 418797 146915 418863 146918
rect 460606 146916 460612 146918
rect 460676 146978 460682 146980
rect 460890 146978 460950 147054
rect 479190 147052 479196 147054
rect 479260 147052 479266 147116
rect 460676 146918 460950 146978
rect 460676 146916 460682 146918
rect 18781 146844 18847 146845
rect 18781 146842 18828 146844
rect 18736 146840 18828 146842
rect 18736 146784 18786 146840
rect 18736 146782 18828 146784
rect 18781 146780 18828 146782
rect 18892 146780 18898 146844
rect 419206 146780 419212 146844
rect 419276 146842 419282 146844
rect 430573 146842 430639 146845
rect 419276 146840 430639 146842
rect 419276 146784 430578 146840
rect 430634 146784 430639 146840
rect 419276 146782 430639 146784
rect 419276 146780 419282 146782
rect 18781 146779 18847 146780
rect 430573 146779 430639 146782
rect 456926 146780 456932 146844
rect 456996 146842 457002 146844
rect 475510 146842 475516 146844
rect 456996 146782 475516 146842
rect 456996 146780 457002 146782
rect 475510 146780 475516 146782
rect 475580 146780 475586 146844
rect 388621 146570 388687 146573
rect 498510 146570 498516 146572
rect 388621 146568 498516 146570
rect 388621 146512 388626 146568
rect 388682 146512 498516 146568
rect 388621 146510 498516 146512
rect 388621 146507 388687 146510
rect 498510 146508 498516 146510
rect 498580 146508 498586 146572
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 551502 136444 551508 136508
rect 551572 136506 551578 136508
rect 551921 136506 551987 136509
rect 551572 136504 551987 136506
rect 551572 136448 551926 136504
rect 551982 136448 551987 136504
rect 551572 136446 551987 136448
rect 551572 136444 551578 136446
rect 551921 136443 551987 136446
rect 151118 135764 151124 135828
rect 151188 135826 151194 135828
rect 151261 135826 151327 135829
rect 151188 135824 151327 135826
rect 151188 135768 151266 135824
rect 151322 135768 151327 135824
rect 151188 135766 151327 135768
rect 151188 135764 151194 135766
rect 151261 135763 151327 135766
rect 158713 129706 158779 129709
rect 558913 129706 558979 129709
rect 156558 129704 158779 129706
rect 156558 129648 158718 129704
rect 158774 129648 158779 129704
rect 156558 129646 158779 129648
rect 156558 129190 156618 129646
rect 158713 129643 158779 129646
rect 556570 129704 558979 129706
rect 556570 129648 558918 129704
rect 558974 129648 558979 129704
rect 556570 129646 558979 129648
rect 556570 129190 556630 129646
rect 558913 129643 558979 129646
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 580257 112779 580323 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 579705 99514 579771 99517
rect 583520 99514 584960 99604
rect 579705 99512 584960 99514
rect 579705 99456 579710 99512
rect 579766 99456 584960 99512
rect 579705 99454 584960 99456
rect 579705 99451 579771 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 16757 86866 16823 86869
rect 19382 86866 20056 86924
rect 16757 86864 20056 86866
rect 417877 86866 417943 86869
rect 419398 86866 420072 86924
rect 417877 86864 420072 86866
rect 16757 86808 16762 86864
rect 16818 86808 19442 86864
rect 16757 86806 19442 86808
rect 417877 86808 417882 86864
rect 417938 86808 419458 86864
rect 417877 86806 419458 86808
rect 16757 86803 16823 86806
rect 417877 86803 417943 86806
rect 580441 86186 580507 86189
rect 583520 86186 584960 86276
rect 580441 86184 584960 86186
rect 580441 86128 580446 86184
rect 580502 86128 584960 86184
rect 580441 86126 584960 86128
rect 580441 86123 580507 86126
rect 583520 86036 584960 86126
rect 17125 85914 17191 85917
rect 19382 85914 20056 85972
rect 17125 85912 20056 85914
rect 417049 85914 417115 85917
rect 419398 85914 420072 85972
rect 417049 85912 420072 85914
rect 17125 85856 17130 85912
rect 17186 85856 19442 85912
rect 17125 85854 19442 85856
rect 417049 85856 417054 85912
rect 417110 85856 419458 85912
rect 417049 85854 419458 85856
rect 17125 85851 17191 85854
rect 417049 85851 417115 85854
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 16941 83738 17007 83741
rect 19382 83738 20056 83796
rect 16941 83736 20056 83738
rect 417969 83738 418035 83741
rect 419398 83738 420072 83796
rect 417969 83736 420072 83738
rect 16941 83680 16946 83736
rect 17002 83680 19442 83736
rect 16941 83678 19442 83680
rect 417969 83680 417974 83736
rect 418030 83680 419458 83736
rect 417969 83678 419458 83680
rect 16941 83675 17007 83678
rect 417969 83675 418035 83678
rect 17585 82922 17651 82925
rect 417417 82922 417483 82925
rect 17585 82920 19810 82922
rect 17585 82864 17590 82920
rect 17646 82864 19810 82920
rect 17585 82862 19810 82864
rect 17585 82859 17651 82862
rect 19750 82844 19810 82862
rect 417417 82920 420010 82922
rect 417417 82864 417422 82920
rect 417478 82864 420010 82920
rect 417417 82862 420010 82864
rect 417417 82859 417483 82862
rect 419950 82844 420010 82862
rect 19750 82784 20056 82844
rect 419950 82784 420072 82844
rect 17493 81018 17559 81021
rect 19382 81018 20056 81076
rect 17493 81016 20056 81018
rect 417233 81018 417299 81021
rect 419398 81018 420072 81076
rect 417233 81016 420072 81018
rect 17493 80960 17498 81016
rect 17554 80960 19442 81016
rect 17493 80958 19442 80960
rect 417233 80960 417238 81016
rect 417294 80960 419458 81016
rect 417233 80958 419458 80960
rect 17493 80955 17559 80958
rect 417233 80955 417299 80958
rect 17861 79930 17927 79933
rect 19382 79930 20056 79988
rect 17861 79928 20056 79930
rect 17861 79872 17866 79928
rect 17922 79872 19442 79928
rect 17861 79870 19442 79872
rect 17861 79867 17927 79870
rect 417918 79868 417924 79932
rect 417988 79930 417994 79932
rect 419398 79930 420072 79988
rect 417988 79928 420072 79930
rect 417988 79870 419458 79928
rect 417988 79868 417994 79870
rect 17769 78162 17835 78165
rect 19382 78162 20056 78220
rect 17769 78160 20056 78162
rect 17769 78104 17774 78160
rect 17830 78104 19442 78160
rect 17769 78102 19442 78104
rect 17769 78099 17835 78102
rect 417734 78100 417740 78164
rect 417804 78162 417810 78164
rect 419398 78162 420072 78220
rect 417804 78160 420072 78162
rect 417804 78102 419458 78160
rect 417804 78100 417810 78102
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 17401 59938 17467 59941
rect 19382 59938 20056 59996
rect 17401 59936 20056 59938
rect 17401 59880 17406 59936
rect 17462 59880 19442 59936
rect 17401 59878 19442 59880
rect 17401 59875 17467 59878
rect 417550 59876 417556 59940
rect 417620 59938 417626 59940
rect 419398 59938 420072 59996
rect 417620 59936 420072 59938
rect 417620 59878 419458 59936
rect 417620 59876 417626 59878
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 17309 58306 17375 58309
rect 19382 58306 20056 58364
rect 17309 58304 20056 58306
rect 417601 58306 417667 58309
rect 419398 58306 420072 58364
rect 417601 58304 420072 58306
rect 17309 58248 17314 58304
rect 17370 58248 19442 58304
rect 17309 58246 19442 58248
rect 417601 58248 417606 58304
rect 417662 58248 419458 58304
rect 417601 58246 419458 58248
rect 17309 58243 17375 58246
rect 417601 58243 417667 58246
rect 19190 57972 19196 58036
rect 19260 58034 19266 58036
rect 19750 58034 20056 58092
rect 19260 58032 20056 58034
rect 416773 58034 416839 58037
rect 419398 58034 420072 58092
rect 416773 58032 420072 58034
rect 19260 57974 19810 58032
rect 416773 57976 416778 58032
rect 416834 57976 419458 58032
rect 416773 57974 419458 57976
rect 19260 57972 19266 57974
rect 416773 57971 416839 57974
rect 53465 49876 53531 49877
rect 60641 49876 60707 49877
rect 456977 49876 457043 49877
rect 458081 49876 458147 49877
rect 478505 49876 478571 49877
rect 53456 49874 53462 49876
rect 53374 49814 53462 49874
rect 53456 49812 53462 49814
rect 53526 49812 53532 49876
rect 60641 49872 60670 49876
rect 60734 49874 60740 49876
rect 60641 49816 60646 49872
rect 60641 49812 60670 49816
rect 60734 49814 60798 49874
rect 456977 49872 456998 49876
rect 457062 49874 457068 49876
rect 456977 49816 456982 49872
rect 60734 49812 60740 49814
rect 456977 49812 456998 49816
rect 457062 49814 457134 49874
rect 457062 49812 457068 49814
rect 458080 49812 458086 49876
rect 458150 49874 458156 49876
rect 478480 49874 478486 49876
rect 458150 49814 458238 49874
rect 478414 49814 478486 49874
rect 478550 49872 478571 49876
rect 478566 49816 478571 49872
rect 458150 49812 458156 49814
rect 478480 49812 478486 49814
rect 478550 49812 478571 49816
rect 53465 49811 53531 49812
rect 60641 49811 60707 49812
rect 456977 49811 457043 49812
rect 458081 49811 458147 49812
rect 478505 49811 478571 49812
rect 480897 49876 480963 49877
rect 480897 49872 480934 49876
rect 480998 49874 481004 49876
rect 480897 49816 480902 49872
rect 480897 49812 480934 49816
rect 480998 49814 481054 49874
rect 480998 49812 481004 49814
rect 480897 49811 480963 49812
rect 91001 49740 91067 49741
rect 95877 49740 95943 49741
rect 473353 49740 473419 49741
rect 90992 49738 90998 49740
rect 90910 49678 90998 49738
rect 90992 49676 90998 49678
rect 91062 49676 91068 49740
rect 95877 49736 95894 49740
rect 95958 49738 95964 49740
rect 473312 49738 473318 49740
rect 95877 49680 95882 49736
rect 95877 49676 95894 49680
rect 95958 49678 96034 49738
rect 473262 49678 473318 49738
rect 473382 49736 473419 49740
rect 473414 49680 473419 49736
rect 95958 49676 95964 49678
rect 473312 49676 473318 49678
rect 473382 49676 473419 49680
rect 91001 49675 91067 49676
rect 95877 49675 95943 49676
rect 473353 49675 473419 49676
rect 488257 49740 488323 49741
rect 495893 49740 495959 49741
rect 503529 49740 503595 49741
rect 488257 49736 488278 49740
rect 488342 49738 488348 49740
rect 495888 49738 495894 49740
rect 488257 49680 488262 49736
rect 488257 49676 488278 49680
rect 488342 49678 488414 49738
rect 495802 49678 495894 49738
rect 488342 49676 488348 49678
rect 495888 49676 495894 49678
rect 495958 49676 495964 49740
rect 503504 49738 503510 49740
rect 503438 49678 503510 49738
rect 503574 49736 503595 49740
rect 503590 49680 503595 49736
rect 503504 49676 503510 49678
rect 503574 49676 503595 49680
rect 488257 49675 488323 49676
rect 495893 49675 495959 49676
rect 503529 49675 503595 49676
rect 48313 49604 48379 49605
rect 50797 49604 50863 49605
rect 53649 49604 53715 49605
rect 56041 49604 56107 49605
rect 58525 49604 58591 49605
rect 80973 49604 81039 49605
rect 83549 49604 83615 49605
rect 86033 49604 86099 49605
rect 48288 49602 48294 49604
rect 48222 49542 48294 49602
rect 48358 49600 48379 49604
rect 50736 49602 50742 49604
rect 48374 49544 48379 49600
rect 48288 49540 48294 49542
rect 48358 49540 48379 49544
rect 50706 49542 50742 49602
rect 50806 49600 50863 49604
rect 53592 49602 53598 49604
rect 50858 49544 50863 49600
rect 50736 49540 50742 49542
rect 50806 49540 50863 49544
rect 53558 49542 53598 49602
rect 53662 49600 53715 49604
rect 53710 49544 53715 49600
rect 53592 49540 53598 49542
rect 53662 49540 53715 49544
rect 56040 49540 56046 49604
rect 56110 49602 56116 49604
rect 58488 49602 58494 49604
rect 56110 49542 56198 49602
rect 58434 49542 58494 49602
rect 58558 49600 58591 49604
rect 80928 49602 80934 49604
rect 58586 49544 58591 49600
rect 56110 49540 56116 49542
rect 58488 49540 58494 49542
rect 58558 49540 58591 49544
rect 80882 49542 80934 49602
rect 80998 49600 81039 49604
rect 83512 49602 83518 49604
rect 81034 49544 81039 49600
rect 80928 49540 80934 49542
rect 80998 49540 81039 49544
rect 83458 49542 83518 49602
rect 83582 49600 83615 49604
rect 85960 49602 85966 49604
rect 83610 49544 83615 49600
rect 83512 49540 83518 49542
rect 83582 49540 83615 49544
rect 85942 49542 85966 49602
rect 85960 49540 85966 49542
rect 86030 49600 86099 49604
rect 86030 49544 86038 49600
rect 86094 49544 86099 49600
rect 86030 49540 86099 49544
rect 48313 49539 48379 49540
rect 50797 49539 50863 49540
rect 53649 49539 53715 49540
rect 56041 49539 56107 49540
rect 58525 49539 58591 49540
rect 80973 49539 81039 49540
rect 83549 49539 83615 49540
rect 86033 49539 86099 49540
rect 88241 49604 88307 49605
rect 98545 49604 98611 49605
rect 103513 49604 103579 49605
rect 105997 49604 106063 49605
rect 88241 49600 88278 49604
rect 88342 49602 88348 49604
rect 98472 49602 98478 49604
rect 88241 49544 88246 49600
rect 88241 49540 88278 49544
rect 88342 49542 88398 49602
rect 98454 49542 98478 49602
rect 88342 49540 88348 49542
rect 98472 49540 98478 49542
rect 98542 49600 98611 49604
rect 98542 49544 98550 49600
rect 98606 49544 98611 49600
rect 98542 49540 98611 49544
rect 103504 49540 103510 49604
rect 103574 49602 103580 49604
rect 105952 49602 105958 49604
rect 103574 49542 103666 49602
rect 105906 49542 105958 49602
rect 106022 49600 106063 49604
rect 106058 49544 106063 49600
rect 103574 49540 103580 49542
rect 105952 49540 105958 49542
rect 106022 49540 106063 49544
rect 120912 49540 120918 49604
rect 120982 49602 120988 49604
rect 389265 49602 389331 49605
rect 120982 49600 389331 49602
rect 120982 49544 389270 49600
rect 389326 49544 389331 49600
rect 120982 49542 389331 49544
rect 120982 49540 120988 49542
rect 88241 49539 88307 49540
rect 98545 49539 98611 49540
rect 103513 49539 103579 49540
rect 105997 49539 106063 49540
rect 389265 49539 389331 49542
rect 410701 49602 410767 49605
rect 493409 49604 493475 49605
rect 498469 49604 498535 49605
rect 500953 49604 501019 49605
rect 490992 49602 490998 49604
rect 410701 49600 490998 49602
rect 410701 49544 410706 49600
rect 410762 49544 490998 49600
rect 410701 49542 490998 49544
rect 410701 49539 410767 49542
rect 490992 49540 490998 49542
rect 491062 49540 491068 49604
rect 493409 49600 493446 49604
rect 493510 49602 493516 49604
rect 493409 49544 493414 49600
rect 493409 49540 493446 49544
rect 493510 49542 493566 49602
rect 498469 49600 498478 49604
rect 498542 49602 498548 49604
rect 500920 49602 500926 49604
rect 498469 49544 498474 49600
rect 493510 49540 493516 49542
rect 498469 49540 498478 49544
rect 498542 49542 498626 49602
rect 500862 49542 500926 49602
rect 500990 49600 501019 49604
rect 501014 49544 501019 49600
rect 498542 49540 498548 49542
rect 500920 49540 500926 49542
rect 500990 49540 501019 49544
rect 493409 49539 493475 49540
rect 498469 49539 498535 49540
rect 500953 49539 501019 49540
rect 505921 49604 505987 49605
rect 508497 49604 508563 49605
rect 510981 49604 511047 49605
rect 513373 49604 513439 49605
rect 515857 49604 515923 49605
rect 520917 49604 520983 49605
rect 525885 49604 525951 49605
rect 505921 49600 505958 49604
rect 506022 49602 506028 49604
rect 505921 49544 505926 49600
rect 505921 49540 505958 49544
rect 506022 49542 506078 49602
rect 508497 49600 508542 49604
rect 508606 49602 508612 49604
rect 508497 49544 508502 49600
rect 506022 49540 506028 49542
rect 508497 49540 508542 49544
rect 508606 49542 508654 49602
rect 510981 49600 510990 49604
rect 511054 49602 511060 49604
rect 510981 49544 510986 49600
rect 508606 49540 508612 49542
rect 510981 49540 510990 49544
rect 511054 49542 511138 49602
rect 513373 49600 513438 49604
rect 513373 49544 513378 49600
rect 513434 49544 513438 49600
rect 511054 49540 511060 49542
rect 513373 49540 513438 49544
rect 513502 49602 513508 49604
rect 513502 49542 513530 49602
rect 515857 49600 515886 49604
rect 515950 49602 515956 49604
rect 520912 49602 520918 49604
rect 515857 49544 515862 49600
rect 513502 49540 513508 49542
rect 515857 49540 515886 49544
rect 515950 49542 516014 49602
rect 520826 49542 520918 49602
rect 515950 49540 515956 49542
rect 520912 49540 520918 49542
rect 520982 49540 520988 49604
rect 525885 49600 525950 49604
rect 525885 49544 525890 49600
rect 525946 49544 525950 49600
rect 525885 49540 525950 49544
rect 526014 49602 526020 49604
rect 526014 49542 526042 49602
rect 526014 49540 526020 49542
rect 505921 49539 505987 49540
rect 508497 49539 508563 49540
rect 510981 49539 511047 49540
rect 513373 49539 513439 49540
rect 515857 49539 515923 49540
rect 520917 49539 520983 49540
rect 525885 49539 525951 49540
rect 113398 49404 113404 49468
rect 113468 49466 113474 49468
rect 161013 49466 161079 49469
rect 113468 49464 161079 49466
rect 113468 49408 161018 49464
rect 161074 49408 161079 49464
rect 113468 49406 161079 49408
rect 113468 49404 113474 49406
rect 161013 49403 161079 49406
rect 407757 49466 407823 49469
rect 485998 49466 486004 49468
rect 407757 49464 486004 49466
rect 407757 49408 407762 49464
rect 407818 49408 486004 49464
rect 407757 49406 486004 49408
rect 407757 49403 407823 49406
rect 485998 49404 486004 49406
rect 486068 49404 486074 49468
rect 408125 49330 408191 49333
rect 483422 49330 483428 49332
rect 408125 49328 483428 49330
rect 408125 49272 408130 49328
rect 408186 49272 483428 49328
rect 408125 49270 483428 49272
rect 408125 49267 408191 49270
rect 483422 49268 483428 49270
rect 483492 49268 483498 49332
rect 418654 49132 418660 49196
rect 418724 49194 418730 49196
rect 460974 49194 460980 49196
rect 418724 49134 460980 49194
rect 418724 49132 418730 49134
rect 460974 49132 460980 49134
rect 461044 49132 461050 49196
rect 459461 49060 459527 49061
rect 419942 48996 419948 49060
rect 420012 49058 420018 49060
rect 459461 49058 459508 49060
rect 420012 49056 459508 49058
rect 420012 49000 459466 49056
rect 420012 48998 459508 49000
rect 420012 48996 420018 48998
rect 459461 48996 459508 48998
rect 459572 48996 459578 49060
rect 459461 48995 459527 48996
rect 36813 48242 36879 48245
rect 43161 48244 43227 48245
rect 37038 48242 37044 48244
rect 36813 48240 37044 48242
rect 36813 48184 36818 48240
rect 36874 48184 37044 48240
rect 36813 48182 37044 48184
rect 36813 48179 36879 48182
rect 37038 48180 37044 48182
rect 37108 48180 37114 48244
rect 43110 48242 43116 48244
rect 43070 48182 43116 48242
rect 43180 48240 43227 48244
rect 43222 48184 43227 48240
rect 43110 48180 43116 48182
rect 43180 48180 43227 48184
rect 43161 48179 43227 48180
rect 44173 48244 44239 48245
rect 45369 48244 45435 48245
rect 44173 48240 44220 48244
rect 44284 48242 44290 48244
rect 45318 48242 45324 48244
rect 44173 48184 44178 48240
rect 44173 48180 44220 48184
rect 44284 48182 44330 48242
rect 45278 48182 45324 48242
rect 45388 48240 45435 48244
rect 45430 48184 45435 48240
rect 44284 48180 44290 48182
rect 45318 48180 45324 48182
rect 45388 48180 45435 48184
rect 44173 48179 44239 48180
rect 45369 48179 45435 48180
rect 46565 48244 46631 48245
rect 47577 48244 47643 48245
rect 48681 48244 48747 48245
rect 46565 48240 46612 48244
rect 46676 48242 46682 48244
rect 47526 48242 47532 48244
rect 46565 48184 46570 48240
rect 46565 48180 46612 48184
rect 46676 48182 46722 48242
rect 47486 48182 47532 48242
rect 47596 48240 47643 48244
rect 48630 48242 48636 48244
rect 47638 48184 47643 48240
rect 46676 48180 46682 48182
rect 47526 48180 47532 48182
rect 47596 48180 47643 48184
rect 48590 48182 48636 48242
rect 48700 48240 48747 48244
rect 48742 48184 48747 48240
rect 48630 48180 48636 48182
rect 48700 48180 48747 48184
rect 46565 48179 46631 48180
rect 47577 48179 47643 48180
rect 48681 48179 48747 48180
rect 49693 48242 49759 48245
rect 50102 48242 50108 48244
rect 49693 48240 50108 48242
rect 49693 48184 49698 48240
rect 49754 48184 50108 48240
rect 49693 48182 50108 48184
rect 49693 48179 49759 48182
rect 50102 48180 50108 48182
rect 50172 48242 50178 48244
rect 50245 48242 50311 48245
rect 51441 48244 51507 48245
rect 52361 48244 52427 48245
rect 54569 48244 54635 48245
rect 55857 48244 55923 48245
rect 51390 48242 51396 48244
rect 50172 48240 50311 48242
rect 50172 48184 50250 48240
rect 50306 48184 50311 48240
rect 50172 48182 50311 48184
rect 51350 48182 51396 48242
rect 51460 48240 51507 48244
rect 52310 48242 52316 48244
rect 51502 48184 51507 48240
rect 50172 48180 50178 48182
rect 50245 48179 50311 48182
rect 51390 48180 51396 48182
rect 51460 48180 51507 48184
rect 52270 48182 52316 48242
rect 52380 48240 52427 48244
rect 54518 48242 54524 48244
rect 52422 48184 52427 48240
rect 52310 48180 52316 48182
rect 52380 48180 52427 48184
rect 54478 48182 54524 48242
rect 54588 48240 54635 48244
rect 55806 48242 55812 48244
rect 54630 48184 54635 48240
rect 54518 48180 54524 48182
rect 54588 48180 54635 48184
rect 55766 48182 55812 48242
rect 55876 48240 55923 48244
rect 55918 48184 55923 48240
rect 55806 48180 55812 48182
rect 55876 48180 55923 48184
rect 51441 48179 51507 48180
rect 52361 48179 52427 48180
rect 54569 48179 54635 48180
rect 55857 48179 55923 48180
rect 57973 48244 58039 48245
rect 59537 48244 59603 48245
rect 61193 48244 61259 48245
rect 57973 48240 58020 48244
rect 58084 48242 58090 48244
rect 59486 48242 59492 48244
rect 57973 48184 57978 48240
rect 57973 48180 58020 48184
rect 58084 48182 58130 48242
rect 59446 48182 59492 48242
rect 59556 48240 59603 48244
rect 61142 48242 61148 48244
rect 59598 48184 59603 48240
rect 58084 48180 58090 48182
rect 59486 48180 59492 48182
rect 59556 48180 59603 48184
rect 61102 48182 61148 48242
rect 61212 48240 61259 48244
rect 61254 48184 61259 48240
rect 61142 48180 61148 48182
rect 61212 48180 61259 48184
rect 57973 48179 58039 48180
rect 59537 48179 59603 48180
rect 61193 48179 61259 48180
rect 61377 48242 61443 48245
rect 61694 48242 61700 48244
rect 61377 48240 61700 48242
rect 61377 48184 61382 48240
rect 61438 48184 61700 48240
rect 61377 48182 61700 48184
rect 61377 48179 61443 48182
rect 61694 48180 61700 48182
rect 61764 48180 61770 48244
rect 62205 48242 62271 48245
rect 62798 48242 62804 48244
rect 62205 48240 62804 48242
rect 62205 48184 62210 48240
rect 62266 48184 62804 48240
rect 62205 48182 62804 48184
rect 62205 48179 62271 48182
rect 62798 48180 62804 48182
rect 62868 48180 62874 48244
rect 63534 48180 63540 48244
rect 63604 48242 63610 48244
rect 63953 48242 64019 48245
rect 63604 48240 64019 48242
rect 63604 48184 63958 48240
rect 64014 48184 64019 48240
rect 63604 48182 64019 48184
rect 63604 48180 63610 48182
rect 63953 48179 64019 48182
rect 65057 48242 65123 48245
rect 65977 48244 66043 48245
rect 65190 48242 65196 48244
rect 65057 48240 65196 48242
rect 65057 48184 65062 48240
rect 65118 48184 65196 48240
rect 65057 48182 65196 48184
rect 65057 48179 65123 48182
rect 65190 48180 65196 48182
rect 65260 48180 65266 48244
rect 65926 48242 65932 48244
rect 65886 48182 65932 48242
rect 65996 48240 66043 48244
rect 66038 48184 66043 48240
rect 65926 48180 65932 48182
rect 65996 48180 66043 48184
rect 65977 48179 66043 48180
rect 66253 48244 66319 48245
rect 67633 48244 67699 48245
rect 68369 48244 68435 48245
rect 66253 48240 66300 48244
rect 66364 48242 66370 48244
rect 67582 48242 67588 48244
rect 66253 48184 66258 48240
rect 66253 48180 66300 48184
rect 66364 48182 66410 48242
rect 67542 48182 67588 48242
rect 67652 48240 67699 48244
rect 68318 48242 68324 48244
rect 67694 48184 67699 48240
rect 66364 48180 66370 48182
rect 67582 48180 67588 48182
rect 67652 48180 67699 48184
rect 68278 48182 68324 48242
rect 68388 48240 68435 48244
rect 68430 48184 68435 48240
rect 68318 48180 68324 48182
rect 68388 48180 68435 48184
rect 66253 48179 66319 48180
rect 67633 48179 67699 48180
rect 68369 48179 68435 48180
rect 68553 48242 68619 48245
rect 69749 48244 69815 48245
rect 68686 48242 68692 48244
rect 68553 48240 68692 48242
rect 68553 48184 68558 48240
rect 68614 48184 68692 48240
rect 68553 48182 68692 48184
rect 68553 48179 68619 48182
rect 68686 48180 68692 48182
rect 68756 48180 68762 48244
rect 69749 48240 69796 48244
rect 69860 48242 69866 48244
rect 69749 48184 69754 48240
rect 69749 48180 69796 48184
rect 69860 48182 69906 48242
rect 69860 48180 69866 48182
rect 70894 48180 70900 48244
rect 70964 48242 70970 48244
rect 71129 48242 71195 48245
rect 70964 48240 71195 48242
rect 70964 48184 71134 48240
rect 71190 48184 71195 48240
rect 70964 48182 71195 48184
rect 70964 48180 70970 48182
rect 69749 48179 69815 48180
rect 71129 48179 71195 48182
rect 71773 48242 71839 48245
rect 73245 48244 73311 48245
rect 72182 48242 72188 48244
rect 71773 48240 72188 48242
rect 71773 48184 71778 48240
rect 71834 48184 72188 48240
rect 71773 48182 72188 48184
rect 71773 48179 71839 48182
rect 72182 48180 72188 48182
rect 72252 48180 72258 48244
rect 73245 48240 73292 48244
rect 73356 48242 73362 48244
rect 73245 48184 73250 48240
rect 73245 48180 73292 48184
rect 73356 48182 73402 48242
rect 73356 48180 73362 48182
rect 73654 48180 73660 48244
rect 73724 48242 73730 48244
rect 73797 48242 73863 48245
rect 73724 48240 73863 48242
rect 73724 48184 73802 48240
rect 73858 48184 73863 48240
rect 73724 48182 73863 48184
rect 73724 48180 73730 48182
rect 73245 48179 73311 48180
rect 73797 48179 73863 48182
rect 74349 48244 74415 48245
rect 76097 48244 76163 48245
rect 74349 48240 74396 48244
rect 74460 48242 74466 48244
rect 76046 48242 76052 48244
rect 74349 48184 74354 48240
rect 74349 48180 74396 48184
rect 74460 48182 74506 48242
rect 76006 48182 76052 48242
rect 76116 48240 76163 48244
rect 76158 48184 76163 48240
rect 74460 48180 74466 48182
rect 76046 48180 76052 48182
rect 76116 48180 76163 48184
rect 74349 48179 74415 48180
rect 76097 48179 76163 48180
rect 76373 48242 76439 48245
rect 78029 48244 78095 48245
rect 78489 48244 78555 48245
rect 93577 48244 93643 48245
rect 100937 48244 101003 48245
rect 76966 48242 76972 48244
rect 76373 48240 76972 48242
rect 76373 48184 76378 48240
rect 76434 48184 76972 48240
rect 76373 48182 76972 48184
rect 76373 48179 76439 48182
rect 76966 48180 76972 48182
rect 77036 48180 77042 48244
rect 78029 48240 78076 48244
rect 78140 48242 78146 48244
rect 78438 48242 78444 48244
rect 78029 48184 78034 48240
rect 78029 48180 78076 48184
rect 78140 48182 78186 48242
rect 78398 48182 78444 48242
rect 78508 48240 78555 48244
rect 93526 48242 93532 48244
rect 78550 48184 78555 48240
rect 78140 48180 78146 48182
rect 78438 48180 78444 48182
rect 78508 48180 78555 48184
rect 93486 48182 93532 48242
rect 93596 48240 93643 48244
rect 100886 48242 100892 48244
rect 93638 48184 93643 48240
rect 93526 48180 93532 48182
rect 93596 48180 93643 48184
rect 100846 48182 100892 48242
rect 100956 48240 101003 48244
rect 100998 48184 101003 48240
rect 100886 48180 100892 48182
rect 100956 48180 101003 48184
rect 108614 48180 108620 48244
rect 108684 48242 108690 48244
rect 108849 48242 108915 48245
rect 108684 48240 108915 48242
rect 108684 48184 108854 48240
rect 108910 48184 108915 48240
rect 108684 48182 108915 48184
rect 108684 48180 108690 48182
rect 78029 48179 78095 48180
rect 78489 48179 78555 48180
rect 93577 48179 93643 48180
rect 100937 48179 101003 48180
rect 108849 48179 108915 48182
rect 111006 48180 111012 48244
rect 111076 48242 111082 48244
rect 111149 48242 111215 48245
rect 115841 48244 115907 48245
rect 118601 48244 118667 48245
rect 125961 48244 126027 48245
rect 115790 48242 115796 48244
rect 111076 48240 111215 48242
rect 111076 48184 111154 48240
rect 111210 48184 111215 48240
rect 111076 48182 111215 48184
rect 115750 48182 115796 48242
rect 115860 48240 115907 48244
rect 118550 48242 118556 48244
rect 115902 48184 115907 48240
rect 111076 48180 111082 48182
rect 111149 48179 111215 48182
rect 115790 48180 115796 48182
rect 115860 48180 115907 48184
rect 118510 48182 118556 48242
rect 118620 48240 118667 48244
rect 125910 48242 125916 48244
rect 118662 48184 118667 48240
rect 118550 48180 118556 48182
rect 118620 48180 118667 48184
rect 125870 48182 125916 48242
rect 125980 48240 126027 48244
rect 126022 48184 126027 48240
rect 125910 48180 125916 48182
rect 125980 48180 126027 48184
rect 115841 48179 115907 48180
rect 118601 48179 118667 48180
rect 125961 48179 126027 48180
rect 436093 48244 436159 48245
rect 437013 48244 437079 48245
rect 438117 48244 438183 48245
rect 439589 48244 439655 48245
rect 443085 48244 443151 48245
rect 444281 48244 444347 48245
rect 436093 48240 436140 48244
rect 436204 48242 436210 48244
rect 436093 48184 436098 48240
rect 436093 48180 436140 48184
rect 436204 48182 436250 48242
rect 437013 48240 437060 48244
rect 437124 48242 437130 48244
rect 437013 48184 437018 48240
rect 436204 48180 436210 48182
rect 437013 48180 437060 48184
rect 437124 48182 437170 48242
rect 438117 48240 438164 48244
rect 438228 48242 438234 48244
rect 438117 48184 438122 48240
rect 437124 48180 437130 48182
rect 438117 48180 438164 48184
rect 438228 48182 438274 48242
rect 439589 48240 439636 48244
rect 439700 48242 439706 48244
rect 439589 48184 439594 48240
rect 438228 48180 438234 48182
rect 439589 48180 439636 48184
rect 439700 48182 439746 48242
rect 443085 48240 443132 48244
rect 443196 48242 443202 48244
rect 444230 48242 444236 48244
rect 443085 48184 443090 48240
rect 439700 48180 439706 48182
rect 443085 48180 443132 48184
rect 443196 48182 443242 48242
rect 444190 48182 444236 48242
rect 444300 48240 444347 48244
rect 444342 48184 444347 48240
rect 443196 48180 443202 48182
rect 444230 48180 444236 48182
rect 444300 48180 444347 48184
rect 436093 48179 436159 48180
rect 437013 48179 437079 48180
rect 438117 48179 438183 48180
rect 439589 48179 439655 48180
rect 443085 48179 443151 48180
rect 444281 48179 444347 48180
rect 448237 48244 448303 48245
rect 450629 48244 450695 48245
rect 453573 48244 453639 48245
rect 454585 48244 454651 48245
rect 448237 48240 448284 48244
rect 448348 48242 448354 48244
rect 448237 48184 448242 48240
rect 448237 48180 448284 48184
rect 448348 48182 448394 48242
rect 450629 48240 450676 48244
rect 450740 48242 450746 48244
rect 450629 48184 450634 48240
rect 448348 48180 448354 48182
rect 450629 48180 450676 48184
rect 450740 48182 450786 48242
rect 453573 48240 453620 48244
rect 453684 48242 453690 48244
rect 454534 48242 454540 48244
rect 453573 48184 453578 48240
rect 450740 48180 450746 48182
rect 453573 48180 453620 48184
rect 453684 48182 453730 48242
rect 454494 48182 454540 48242
rect 454604 48240 454651 48244
rect 454646 48184 454651 48240
rect 453684 48180 453690 48182
rect 454534 48180 454540 48182
rect 454604 48180 454651 48184
rect 455638 48180 455644 48244
rect 455708 48242 455714 48244
rect 455873 48242 455939 48245
rect 455708 48240 455939 48242
rect 455708 48184 455878 48240
rect 455934 48184 455939 48240
rect 455708 48182 455939 48184
rect 455708 48180 455714 48182
rect 448237 48179 448303 48180
rect 450629 48179 450695 48180
rect 453573 48179 453639 48180
rect 454585 48179 454651 48180
rect 455873 48179 455939 48182
rect 458357 48244 458423 48245
rect 461669 48244 461735 48245
rect 462773 48244 462839 48245
rect 463509 48244 463575 48245
rect 463877 48244 463943 48245
rect 465165 48244 465231 48245
rect 465901 48244 465967 48245
rect 466269 48244 466335 48245
rect 467557 48244 467623 48245
rect 468293 48244 468359 48245
rect 468661 48244 468727 48245
rect 458357 48240 458404 48244
rect 458468 48242 458474 48244
rect 458357 48184 458362 48240
rect 458357 48180 458404 48184
rect 458468 48182 458514 48242
rect 461669 48240 461716 48244
rect 461780 48242 461786 48244
rect 461669 48184 461674 48240
rect 458468 48180 458474 48182
rect 461669 48180 461716 48184
rect 461780 48182 461826 48242
rect 462773 48240 462820 48244
rect 462884 48242 462890 48244
rect 462773 48184 462778 48240
rect 461780 48180 461786 48182
rect 462773 48180 462820 48184
rect 462884 48182 462930 48242
rect 463509 48240 463556 48244
rect 463620 48242 463626 48244
rect 463509 48184 463514 48240
rect 462884 48180 462890 48182
rect 463509 48180 463556 48184
rect 463620 48182 463666 48242
rect 463877 48240 463924 48244
rect 463988 48242 463994 48244
rect 463877 48184 463882 48240
rect 463620 48180 463626 48182
rect 463877 48180 463924 48184
rect 463988 48182 464034 48242
rect 465165 48240 465212 48244
rect 465276 48242 465282 48244
rect 465165 48184 465170 48240
rect 463988 48180 463994 48182
rect 465165 48180 465212 48184
rect 465276 48182 465322 48242
rect 465901 48240 465948 48244
rect 466012 48242 466018 48244
rect 465901 48184 465906 48240
rect 465276 48180 465282 48182
rect 465901 48180 465948 48184
rect 466012 48182 466058 48242
rect 466269 48240 466316 48244
rect 466380 48242 466386 48244
rect 466269 48184 466274 48240
rect 466012 48180 466018 48182
rect 466269 48180 466316 48184
rect 466380 48182 466426 48242
rect 467557 48240 467604 48244
rect 467668 48242 467674 48244
rect 467557 48184 467562 48240
rect 466380 48180 466386 48182
rect 467557 48180 467604 48184
rect 467668 48182 467714 48242
rect 468293 48240 468340 48244
rect 468404 48242 468410 48244
rect 468293 48184 468298 48240
rect 467668 48180 467674 48182
rect 468293 48180 468340 48184
rect 468404 48182 468450 48242
rect 468661 48240 468708 48244
rect 468772 48242 468778 48244
rect 469213 48242 469279 48245
rect 470869 48244 470935 48245
rect 471237 48244 471303 48245
rect 472157 48244 472223 48245
rect 474365 48244 474431 48245
rect 475653 48244 475719 48245
rect 476941 48244 477007 48245
rect 478045 48244 478111 48245
rect 469806 48242 469812 48244
rect 468661 48184 468666 48240
rect 468404 48180 468410 48182
rect 468661 48180 468708 48184
rect 468772 48182 468818 48242
rect 469213 48240 469812 48242
rect 469213 48184 469218 48240
rect 469274 48184 469812 48240
rect 469213 48182 469812 48184
rect 468772 48180 468778 48182
rect 458357 48179 458423 48180
rect 461669 48179 461735 48180
rect 462773 48179 462839 48180
rect 463509 48179 463575 48180
rect 463877 48179 463943 48180
rect 465165 48179 465231 48180
rect 465901 48179 465967 48180
rect 466269 48179 466335 48180
rect 467557 48179 467623 48180
rect 468293 48179 468359 48180
rect 468661 48179 468727 48180
rect 469213 48179 469279 48182
rect 469806 48180 469812 48182
rect 469876 48180 469882 48244
rect 470869 48240 470916 48244
rect 470980 48242 470986 48244
rect 470869 48184 470874 48240
rect 470869 48180 470916 48184
rect 470980 48182 471026 48242
rect 471237 48240 471284 48244
rect 471348 48242 471354 48244
rect 471237 48184 471242 48240
rect 470980 48180 470986 48182
rect 471237 48180 471284 48184
rect 471348 48182 471394 48242
rect 472157 48240 472204 48244
rect 472268 48242 472274 48244
rect 472157 48184 472162 48240
rect 471348 48180 471354 48182
rect 472157 48180 472204 48184
rect 472268 48182 472314 48242
rect 474365 48240 474412 48244
rect 474476 48242 474482 48244
rect 474365 48184 474370 48240
rect 472268 48180 472274 48182
rect 474365 48180 474412 48184
rect 474476 48182 474522 48242
rect 475653 48240 475700 48244
rect 475764 48242 475770 48244
rect 475653 48184 475658 48240
rect 474476 48180 474482 48182
rect 475653 48180 475700 48184
rect 475764 48182 475810 48242
rect 476941 48240 476988 48244
rect 477052 48242 477058 48244
rect 476941 48184 476946 48240
rect 475764 48180 475770 48182
rect 476941 48180 476988 48184
rect 477052 48182 477098 48242
rect 478045 48240 478092 48244
rect 478156 48242 478162 48244
rect 478045 48184 478050 48240
rect 477052 48180 477058 48182
rect 478045 48180 478092 48184
rect 478156 48182 478202 48242
rect 478156 48180 478162 48182
rect 470869 48179 470935 48180
rect 471237 48179 471303 48180
rect 472157 48179 472223 48180
rect 474365 48179 474431 48180
rect 475653 48179 475719 48180
rect 476941 48179 477007 48180
rect 478045 48179 478111 48180
rect 19517 48106 19583 48109
rect 63861 48108 63927 48109
rect 71037 48108 71103 48109
rect 445293 48108 445359 48109
rect 446397 48108 446463 48109
rect 40534 48106 40540 48108
rect 19517 48104 40540 48106
rect 19517 48048 19522 48104
rect 19578 48048 40540 48104
rect 19517 48046 40540 48048
rect 19517 48043 19583 48046
rect 40534 48044 40540 48046
rect 40604 48044 40610 48108
rect 41822 48044 41828 48108
rect 41892 48044 41898 48108
rect 63861 48104 63908 48108
rect 63972 48106 63978 48108
rect 63861 48048 63866 48104
rect 63861 48044 63908 48048
rect 63972 48046 64018 48106
rect 71037 48104 71084 48108
rect 71148 48106 71154 48108
rect 71037 48048 71042 48104
rect 63972 48044 63978 48046
rect 71037 48044 71084 48048
rect 71148 48046 71194 48106
rect 71148 48044 71154 48046
rect 123334 48044 123340 48108
rect 123404 48106 123410 48108
rect 389214 48106 389220 48108
rect 123404 48046 389220 48106
rect 123404 48044 123410 48046
rect 389214 48044 389220 48046
rect 389284 48044 389290 48108
rect 419390 48044 419396 48108
rect 419460 48106 419466 48108
rect 440550 48106 440556 48108
rect 419460 48046 440556 48106
rect 419460 48044 419466 48046
rect 440550 48044 440556 48046
rect 440620 48044 440626 48108
rect 445293 48104 445340 48108
rect 445404 48106 445410 48108
rect 445293 48048 445298 48104
rect 445293 48044 445340 48048
rect 445404 48046 445450 48106
rect 446397 48104 446444 48108
rect 446508 48106 446514 48108
rect 446397 48048 446402 48104
rect 445404 48044 445410 48046
rect 446397 48044 446444 48048
rect 446508 48046 446554 48106
rect 446508 48044 446514 48046
rect 448646 48044 448652 48108
rect 448716 48106 448722 48108
rect 449525 48106 449591 48109
rect 448716 48104 449591 48106
rect 448716 48048 449530 48104
rect 449586 48048 449591 48104
rect 448716 48046 449591 48048
rect 448716 48044 448722 48046
rect 18781 47970 18847 47973
rect 39614 47970 39620 47972
rect 18781 47968 39620 47970
rect 18781 47912 18786 47968
rect 18842 47912 39620 47968
rect 18781 47910 39620 47912
rect 18781 47907 18847 47910
rect 39614 47908 39620 47910
rect 39684 47908 39690 47972
rect 18689 47834 18755 47837
rect 38510 47834 38516 47836
rect 18689 47832 38516 47834
rect 18689 47776 18694 47832
rect 18750 47776 38516 47832
rect 18689 47774 38516 47776
rect 18689 47771 18755 47774
rect 38510 47772 38516 47774
rect 38580 47772 38586 47836
rect 18638 47636 18644 47700
rect 18708 47698 18714 47700
rect 41830 47698 41890 48044
rect 63861 48043 63927 48044
rect 71037 48043 71103 48044
rect 445293 48043 445359 48044
rect 446397 48043 446463 48044
rect 449525 48043 449591 48046
rect 452285 48108 452351 48109
rect 452285 48104 452332 48108
rect 452396 48106 452402 48108
rect 452285 48048 452290 48104
rect 452285 48044 452332 48048
rect 452396 48046 452442 48106
rect 452396 48044 452402 48046
rect 453430 48044 453436 48108
rect 453500 48106 453506 48108
rect 453941 48106 454007 48109
rect 453500 48104 454007 48106
rect 453500 48048 453946 48104
rect 454002 48048 454007 48104
rect 453500 48046 454007 48048
rect 453500 48044 453506 48046
rect 452285 48043 452351 48044
rect 453941 48043 454007 48046
rect 456977 48106 457043 48109
rect 469121 48106 469187 48109
rect 456977 48104 469187 48106
rect 456977 48048 456982 48104
rect 457038 48048 469126 48104
rect 469182 48048 469187 48104
rect 456977 48046 469187 48048
rect 456977 48043 457043 48046
rect 469121 48043 469187 48046
rect 60641 47970 60707 47973
rect 79174 47970 79180 47972
rect 60641 47968 79180 47970
rect 60641 47912 60646 47968
rect 60702 47912 79180 47968
rect 60641 47910 79180 47912
rect 60641 47907 60707 47910
rect 79174 47908 79180 47910
rect 79244 47908 79250 47972
rect 404997 47970 405063 47973
rect 475878 47970 475884 47972
rect 404997 47968 475884 47970
rect 404997 47912 405002 47968
rect 405058 47912 475884 47968
rect 404997 47910 475884 47912
rect 404997 47907 405063 47910
rect 475878 47908 475884 47910
rect 475948 47908 475954 47972
rect 405181 47834 405247 47837
rect 473302 47834 473308 47836
rect 405181 47832 473308 47834
rect 405181 47776 405186 47832
rect 405242 47776 473308 47832
rect 405181 47774 473308 47776
rect 405181 47771 405247 47774
rect 473302 47772 473308 47774
rect 473372 47772 473378 47836
rect 18708 47638 41890 47698
rect 18708 47636 18714 47638
rect 415894 47636 415900 47700
rect 415964 47698 415970 47700
rect 455822 47698 455828 47700
rect 415964 47638 455828 47698
rect 415964 47636 415970 47638
rect 455822 47636 455828 47638
rect 455892 47636 455898 47700
rect 459921 47698 459987 47701
rect 460606 47698 460612 47700
rect 459921 47696 460612 47698
rect 459921 47640 459926 47696
rect 459982 47640 460612 47696
rect 459921 47638 460612 47640
rect 459921 47635 459987 47638
rect 460606 47636 460612 47638
rect 460676 47698 460682 47700
rect 479190 47698 479196 47700
rect 460676 47638 479196 47698
rect 460676 47636 460682 47638
rect 479190 47636 479196 47638
rect 479260 47636 479266 47700
rect 18965 47562 19031 47565
rect 57053 47564 57119 47565
rect 447501 47564 447567 47565
rect 35934 47562 35940 47564
rect 18965 47560 35940 47562
rect 18965 47504 18970 47560
rect 19026 47504 35940 47560
rect 18965 47502 35940 47504
rect 18965 47499 19031 47502
rect 35934 47500 35940 47502
rect 36004 47500 36010 47564
rect 57053 47562 57100 47564
rect 56972 47560 57100 47562
rect 57164 47562 57170 47564
rect 75678 47562 75684 47564
rect 56972 47504 57058 47560
rect 56972 47502 57100 47504
rect 57053 47500 57100 47502
rect 57164 47502 75684 47562
rect 57164 47500 57170 47502
rect 75678 47500 75684 47502
rect 75748 47500 75754 47564
rect 419206 47500 419212 47564
rect 419276 47562 419282 47564
rect 447501 47562 447548 47564
rect 419276 47502 431970 47562
rect 447456 47560 447548 47562
rect 447456 47504 447506 47560
rect 447456 47502 447548 47504
rect 419276 47500 419282 47502
rect 57053 47499 57119 47500
rect 431910 47426 431970 47502
rect 447501 47500 447548 47502
rect 447612 47500 447618 47564
rect 447501 47499 447567 47500
rect 450077 47428 450143 47429
rect 442022 47426 442028 47428
rect 431910 47366 442028 47426
rect 442022 47364 442028 47366
rect 442092 47364 442098 47428
rect 450077 47426 450124 47428
rect 449996 47424 450124 47426
rect 450188 47426 450194 47428
rect 450445 47426 450511 47429
rect 451273 47428 451339 47429
rect 450188 47424 450511 47426
rect 449996 47368 450082 47424
rect 450188 47368 450450 47424
rect 450506 47368 450511 47424
rect 449996 47366 450124 47368
rect 450077 47364 450124 47366
rect 450188 47366 450511 47368
rect 450188 47364 450194 47366
rect 450077 47363 450143 47364
rect 450445 47363 450511 47366
rect 451222 47364 451228 47428
rect 451292 47426 451339 47428
rect 451292 47424 451384 47426
rect 451334 47368 451384 47424
rect 451292 47366 451384 47368
rect 451292 47364 451339 47366
rect 451273 47363 451339 47364
rect 416221 47290 416287 47293
rect 523350 47290 523356 47292
rect 416221 47288 523356 47290
rect 416221 47232 416226 47288
rect 416282 47232 523356 47288
rect 416221 47230 523356 47232
rect 416221 47227 416287 47230
rect 523350 47228 523356 47230
rect 523420 47228 523426 47292
rect 416405 47154 416471 47157
rect 518382 47154 518388 47156
rect 416405 47152 518388 47154
rect 416405 47096 416410 47152
rect 416466 47096 518388 47152
rect 416405 47094 518388 47096
rect 416405 47091 416471 47094
rect 518382 47092 518388 47094
rect 518452 47092 518458 47156
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 193806 31724 193812 31788
rect 193876 31786 193882 31788
rect 583526 31786 583586 32950
rect 193876 31726 583586 31786
rect 193876 31724 193882 31726
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 193990 19348 193996 19412
rect 194060 19410 194066 19412
rect 583526 19410 583586 19622
rect 194060 19350 583586 19410
rect 194060 19348 194066 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 193812 682076 193876 682140
rect 186268 681940 186332 682004
rect 193996 681804 194060 681868
rect 186268 678132 186332 678196
rect 550956 585168 551020 585172
rect 550956 585112 551006 585168
rect 551006 585112 551020 585168
rect 550956 585108 551020 585112
rect 441660 498128 441724 498132
rect 441660 498072 441674 498128
rect 441674 498072 441724 498128
rect 441660 498068 441724 498072
rect 445340 498068 445404 498132
rect 448652 498068 448716 498132
rect 452332 498068 452396 498132
rect 456196 498068 456260 498132
rect 473492 498068 473556 498132
rect 480852 498068 480916 498132
rect 486004 497932 486068 497996
rect 453436 497524 453500 497588
rect 437060 497252 437124 497316
rect 436140 497176 436204 497180
rect 436140 497120 436154 497176
rect 436154 497120 436204 497176
rect 436140 497116 436204 497120
rect 455828 497116 455892 497180
rect 483428 497116 483492 497180
rect 444236 496980 444300 497044
rect 448284 496980 448348 497044
rect 450676 496980 450740 497044
rect 456932 497040 456996 497044
rect 456932 496984 456946 497040
rect 456946 496984 456996 497040
rect 456932 496980 456996 496984
rect 459324 496980 459388 497044
rect 460612 496980 460676 497044
rect 470916 496980 470980 497044
rect 476068 497040 476132 497044
rect 476068 496984 476118 497040
rect 476118 496984 476132 497040
rect 476068 496980 476132 496984
rect 438348 496844 438412 496908
rect 439636 496844 439700 496908
rect 440556 496844 440620 496908
rect 443132 496904 443196 496908
rect 443132 496848 443146 496904
rect 443146 496848 443196 496904
rect 443132 496844 443196 496848
rect 446444 496844 446508 496908
rect 447548 496844 447612 496908
rect 449940 496904 450004 496908
rect 449940 496848 449954 496904
rect 449954 496848 450004 496904
rect 449940 496844 450004 496848
rect 451044 496844 451108 496908
rect 453620 496844 453684 496908
rect 454540 496844 454604 496908
rect 458036 496844 458100 496908
rect 458404 496844 458468 496908
rect 460980 496904 461044 496908
rect 460980 496848 460994 496904
rect 460994 496848 461044 496904
rect 460980 496844 461044 496848
rect 463556 496844 463620 496908
rect 465948 496844 466012 496908
rect 468340 496844 468404 496908
rect 478460 496844 478524 496908
rect 3372 466516 3436 466580
rect 193996 462844 194060 462908
rect 418660 462708 418724 462772
rect 193812 457404 193876 457468
rect 19196 455636 19260 455700
rect 418108 454548 418172 454612
rect 19012 453324 19076 453388
rect 192340 453052 192404 453116
rect 191604 452644 191668 452708
rect 418844 450468 418908 450532
rect 193996 450332 194060 450396
rect 415900 450196 415964 450260
rect 389220 449652 389284 449716
rect 193812 449244 193876 449308
rect 150940 435236 151004 435300
rect 550838 433468 550902 433532
rect 417924 359892 417988 359956
rect 90998 349888 91062 349892
rect 90998 349832 91006 349888
rect 91006 349832 91062 349888
rect 90998 349828 91062 349832
rect 93446 349888 93510 349892
rect 93446 349832 93490 349888
rect 93490 349832 93510 349888
rect 93446 349828 93510 349832
rect 98478 349828 98542 349892
rect 103510 349888 103574 349892
rect 103510 349832 103518 349888
rect 103518 349832 103574 349888
rect 103510 349828 103574 349832
rect 478486 349888 478550 349892
rect 478486 349832 478510 349888
rect 478510 349832 478550 349888
rect 478486 349828 478550 349832
rect 483518 349888 483582 349892
rect 483518 349832 483534 349888
rect 483534 349832 483582 349888
rect 483518 349828 483582 349832
rect 485966 349888 486030 349892
rect 485966 349832 486018 349888
rect 486018 349832 486030 349888
rect 485966 349828 486030 349832
rect 495894 349828 495958 349892
rect 452374 349692 452438 349756
rect 488278 349752 488342 349756
rect 488278 349696 488318 349752
rect 488318 349696 488342 349752
rect 488278 349692 488342 349696
rect 490998 349752 491062 349756
rect 490998 349696 491022 349752
rect 491022 349696 491062 349752
rect 490998 349692 491062 349696
rect 508542 349752 508606 349756
rect 508542 349696 508558 349752
rect 508558 349696 508606 349752
rect 508542 349692 508606 349696
rect 520918 349752 520982 349756
rect 520918 349696 520922 349752
rect 520922 349696 520978 349752
rect 520978 349696 520982 349752
rect 520918 349692 520982 349696
rect 38230 349556 38294 349620
rect 50742 349616 50806 349620
rect 50742 349560 50802 349616
rect 50802 349560 50806 349616
rect 50742 349556 50806 349560
rect 56046 349616 56110 349620
rect 56046 349560 56102 349616
rect 56102 349560 56110 349616
rect 56046 349556 56110 349560
rect 58494 349616 58558 349620
rect 58494 349560 58530 349616
rect 58530 349560 58558 349616
rect 58494 349556 58558 349560
rect 61078 349616 61142 349620
rect 61078 349560 61106 349616
rect 61106 349560 61142 349616
rect 61078 349556 61142 349560
rect 62846 349616 62910 349620
rect 62846 349560 62854 349616
rect 62854 349560 62910 349616
rect 62846 349556 62910 349560
rect 68694 349616 68758 349620
rect 68694 349560 68742 349616
rect 68742 349560 68758 349616
rect 68694 349556 68758 349560
rect 72230 349616 72294 349620
rect 72230 349560 72238 349616
rect 72238 349560 72294 349616
rect 72230 349556 72294 349560
rect 505958 349616 506022 349620
rect 505958 349560 505982 349616
rect 505982 349560 506022 349616
rect 505958 349556 506022 349560
rect 515886 349616 515950 349620
rect 515886 349560 515918 349616
rect 515918 349560 515950 349616
rect 515886 349556 515950 349560
rect 480852 349148 480916 349212
rect 53604 349072 53668 349076
rect 53604 349016 53654 349072
rect 53654 349016 53668 349072
rect 53604 349012 53668 349016
rect 61884 349012 61948 349076
rect 68324 349072 68388 349076
rect 68324 349016 68374 349072
rect 68374 349016 68388 349072
rect 68324 349012 68388 349016
rect 78444 349072 78508 349076
rect 78444 349016 78494 349072
rect 78494 349016 78508 349072
rect 78444 349012 78508 349016
rect 85988 349072 86052 349076
rect 85988 349016 86038 349072
rect 86038 349016 86052 349072
rect 85988 349012 86052 349016
rect 88196 349012 88260 349076
rect 498516 349072 498580 349076
rect 498516 349016 498530 349072
rect 498530 349016 498580 349072
rect 498516 349012 498580 349016
rect 500908 349072 500972 349076
rect 500908 349016 500958 349072
rect 500958 349016 500972 349072
rect 500908 349012 500972 349016
rect 503484 349072 503548 349076
rect 503484 349016 503498 349072
rect 503498 349016 503548 349072
rect 503484 349012 503548 349016
rect 511028 349072 511092 349076
rect 511028 349016 511042 349072
rect 511042 349016 511092 349072
rect 511028 349012 511092 349016
rect 523356 349072 523420 349076
rect 523356 349016 523370 349072
rect 523370 349016 523420 349072
rect 523356 349012 523420 349016
rect 74396 348528 74460 348532
rect 74396 348472 74410 348528
rect 74410 348472 74460 348528
rect 74396 348468 74460 348472
rect 419764 347788 419828 347852
rect 36124 347712 36188 347716
rect 36124 347656 36174 347712
rect 36174 347656 36188 347712
rect 36124 347652 36188 347656
rect 39620 347712 39684 347716
rect 39620 347656 39634 347712
rect 39634 347656 39684 347712
rect 39620 347652 39684 347656
rect 43116 347652 43180 347716
rect 44220 347712 44284 347716
rect 44220 347656 44234 347712
rect 44234 347656 44284 347712
rect 44220 347652 44284 347656
rect 45324 347712 45388 347716
rect 45324 347656 45374 347712
rect 45374 347656 45388 347712
rect 45324 347652 45388 347656
rect 46612 347712 46676 347716
rect 46612 347656 46626 347712
rect 46626 347656 46676 347712
rect 46612 347652 46676 347656
rect 47532 347712 47596 347716
rect 47532 347656 47582 347712
rect 47582 347656 47596 347712
rect 47532 347652 47596 347656
rect 48636 347712 48700 347716
rect 48636 347656 48650 347712
rect 48650 347656 48700 347712
rect 48636 347652 48700 347656
rect 50108 347712 50172 347716
rect 50108 347656 50122 347712
rect 50122 347656 50172 347712
rect 50108 347652 50172 347656
rect 51212 347712 51276 347716
rect 51212 347656 51262 347712
rect 51262 347656 51276 347712
rect 51212 347652 51276 347656
rect 52316 347712 52380 347716
rect 52316 347656 52366 347712
rect 52366 347656 52380 347712
rect 52316 347652 52380 347656
rect 53420 347712 53484 347716
rect 53420 347656 53470 347712
rect 53470 347656 53484 347712
rect 53420 347652 53484 347656
rect 63540 347652 63604 347716
rect 63908 347652 63972 347716
rect 65196 347712 65260 347716
rect 65196 347656 65210 347712
rect 65210 347656 65260 347712
rect 65196 347652 65260 347656
rect 65932 347712 65996 347716
rect 65932 347656 65982 347712
rect 65982 347656 65996 347712
rect 65932 347652 65996 347656
rect 66300 347712 66364 347716
rect 66300 347656 66314 347712
rect 66314 347656 66364 347712
rect 66300 347652 66364 347656
rect 67588 347652 67652 347716
rect 71268 347652 71332 347716
rect 73292 347712 73356 347716
rect 73292 347656 73306 347712
rect 73306 347656 73356 347712
rect 73292 347652 73356 347656
rect 73660 347712 73724 347716
rect 73660 347656 73710 347712
rect 73710 347656 73724 347712
rect 73660 347652 73724 347656
rect 75684 347652 75748 347716
rect 76052 347712 76116 347716
rect 76052 347656 76102 347712
rect 76102 347656 76116 347712
rect 76052 347652 76116 347656
rect 76972 347652 77036 347716
rect 78076 347712 78140 347716
rect 78076 347656 78090 347712
rect 78090 347656 78140 347712
rect 78076 347652 78140 347656
rect 79180 347712 79244 347716
rect 79180 347656 79194 347712
rect 79194 347656 79244 347712
rect 79180 347652 79244 347656
rect 81020 347712 81084 347716
rect 81020 347656 81070 347712
rect 81070 347656 81084 347712
rect 81020 347652 81084 347656
rect 83596 347712 83660 347716
rect 83596 347656 83646 347712
rect 83646 347656 83660 347712
rect 83596 347652 83660 347656
rect 95924 347652 95988 347716
rect 100892 347712 100956 347716
rect 100892 347656 100942 347712
rect 100942 347656 100956 347712
rect 100892 347652 100956 347656
rect 106044 347712 106108 347716
rect 106044 347656 106094 347712
rect 106094 347656 106108 347712
rect 106044 347652 106108 347656
rect 108620 347712 108684 347716
rect 108620 347656 108670 347712
rect 108670 347656 108684 347712
rect 108620 347652 108684 347656
rect 111012 347712 111076 347716
rect 111012 347656 111062 347712
rect 111062 347656 111076 347712
rect 111012 347652 111076 347656
rect 113404 347712 113468 347716
rect 113404 347656 113454 347712
rect 113454 347656 113468 347712
rect 113404 347652 113468 347656
rect 115796 347712 115860 347716
rect 115796 347656 115846 347712
rect 115846 347656 115860 347712
rect 115796 347652 115860 347656
rect 118556 347712 118620 347716
rect 118556 347656 118606 347712
rect 118606 347656 118620 347712
rect 118556 347652 118620 347656
rect 120948 347712 121012 347716
rect 120948 347656 120998 347712
rect 120998 347656 121012 347712
rect 120948 347652 121012 347656
rect 123340 347712 123404 347716
rect 123340 347656 123390 347712
rect 123390 347656 123404 347712
rect 123340 347652 123404 347656
rect 125916 347712 125980 347716
rect 125916 347656 125966 347712
rect 125966 347656 125980 347712
rect 125916 347652 125980 347656
rect 48268 347516 48332 347580
rect 436140 347712 436204 347716
rect 436140 347656 436154 347712
rect 436154 347656 436204 347712
rect 436140 347652 436204 347656
rect 437060 347712 437124 347716
rect 437060 347656 437074 347712
rect 437074 347656 437124 347712
rect 437060 347652 437124 347656
rect 438164 347652 438228 347716
rect 439636 347712 439700 347716
rect 439636 347656 439650 347712
rect 439650 347656 439700 347712
rect 439636 347652 439700 347656
rect 440556 347712 440620 347716
rect 440556 347656 440570 347712
rect 440570 347656 440620 347712
rect 440556 347652 440620 347656
rect 441660 347712 441724 347716
rect 441660 347656 441674 347712
rect 441674 347656 441724 347712
rect 441660 347652 441724 347656
rect 443132 347712 443196 347716
rect 443132 347656 443146 347712
rect 443146 347656 443196 347712
rect 443132 347652 443196 347656
rect 444236 347712 444300 347716
rect 444236 347656 444250 347712
rect 444250 347656 444300 347712
rect 444236 347652 444300 347656
rect 445340 347712 445404 347716
rect 445340 347656 445354 347712
rect 445354 347656 445404 347712
rect 445340 347652 445404 347656
rect 446444 347712 446508 347716
rect 446444 347656 446458 347712
rect 446458 347656 446508 347712
rect 446444 347652 446508 347656
rect 447548 347652 447612 347716
rect 448284 347712 448348 347716
rect 448284 347656 448298 347712
rect 448298 347656 448348 347712
rect 448284 347652 448348 347656
rect 448652 347652 448716 347716
rect 450124 347652 450188 347716
rect 450676 347712 450740 347716
rect 450676 347656 450690 347712
rect 450690 347656 450740 347712
rect 450676 347652 450740 347656
rect 451412 347712 451476 347716
rect 451412 347656 451426 347712
rect 451426 347656 451476 347712
rect 451412 347652 451476 347656
rect 453436 347652 453500 347716
rect 453620 347712 453684 347716
rect 453620 347656 453634 347712
rect 453634 347656 453684 347712
rect 453620 347652 453684 347656
rect 454540 347652 454604 347716
rect 455828 347712 455892 347716
rect 455828 347656 455842 347712
rect 455842 347656 455892 347712
rect 455828 347652 455892 347656
rect 456196 347712 456260 347716
rect 456196 347656 456210 347712
rect 456210 347656 456260 347712
rect 456196 347652 456260 347656
rect 456932 347712 456996 347716
rect 456932 347656 456982 347712
rect 456982 347656 456996 347712
rect 456932 347652 456996 347656
rect 458036 347712 458100 347716
rect 458036 347656 458086 347712
rect 458086 347656 458100 347712
rect 458036 347652 458100 347656
rect 458404 347712 458468 347716
rect 458404 347656 458418 347712
rect 458418 347656 458468 347712
rect 458404 347652 458468 347656
rect 459508 347712 459572 347716
rect 459508 347656 459522 347712
rect 459522 347656 459572 347712
rect 459508 347652 459572 347656
rect 460980 347712 461044 347716
rect 460980 347656 460994 347712
rect 460994 347656 461044 347712
rect 460980 347652 461044 347656
rect 461716 347652 461780 347716
rect 462820 347712 462884 347716
rect 462820 347656 462834 347712
rect 462834 347656 462884 347712
rect 462820 347652 462884 347656
rect 463556 347712 463620 347716
rect 463556 347656 463570 347712
rect 463570 347656 463620 347712
rect 463556 347652 463620 347656
rect 463924 347712 463988 347716
rect 463924 347656 463938 347712
rect 463938 347656 463988 347712
rect 463924 347652 463988 347656
rect 465212 347712 465276 347716
rect 465212 347656 465226 347712
rect 465226 347656 465276 347712
rect 465212 347652 465276 347656
rect 466316 347652 466380 347716
rect 467604 347652 467668 347716
rect 468340 347516 468404 347580
rect 468708 347712 468772 347716
rect 468708 347656 468722 347712
rect 468722 347656 468772 347712
rect 468708 347652 468772 347656
rect 469812 347712 469876 347716
rect 469812 347656 469826 347712
rect 469826 347656 469876 347712
rect 469812 347652 469876 347656
rect 471284 347712 471348 347716
rect 471284 347656 471298 347712
rect 471298 347656 471348 347712
rect 471284 347652 471348 347656
rect 472204 347652 472268 347716
rect 473308 347712 473372 347716
rect 473308 347656 473358 347712
rect 473358 347656 473372 347712
rect 473308 347652 473372 347656
rect 474412 347712 474476 347716
rect 474412 347656 474426 347712
rect 474426 347656 474476 347712
rect 474412 347652 474476 347656
rect 475700 347712 475764 347716
rect 475700 347656 475714 347712
rect 475714 347656 475764 347712
rect 475700 347652 475764 347656
rect 476988 347712 477052 347716
rect 476988 347656 477002 347712
rect 477002 347656 477052 347712
rect 476988 347652 477052 347656
rect 478092 347712 478156 347716
rect 478092 347656 478106 347712
rect 478106 347656 478156 347712
rect 478092 347652 478156 347656
rect 479196 347712 479260 347716
rect 479196 347656 479210 347712
rect 479210 347656 479260 347712
rect 479196 347652 479260 347656
rect 513420 347712 513484 347716
rect 513420 347656 513434 347712
rect 513434 347656 513484 347712
rect 513420 347652 513484 347656
rect 518388 347712 518452 347716
rect 518388 347656 518402 347712
rect 518402 347656 518452 347712
rect 518388 347652 518452 347656
rect 525932 347712 525996 347716
rect 525932 347656 525946 347712
rect 525946 347656 525996 347712
rect 525932 347652 525996 347656
rect 470364 347516 470428 347580
rect 55812 347380 55876 347444
rect 58204 347380 58268 347444
rect 59492 347380 59556 347444
rect 70900 347380 70964 347444
rect 473492 347380 473556 347444
rect 37228 347304 37292 347308
rect 37228 347248 37242 347304
rect 37242 347248 37292 347304
rect 37228 347244 37292 347248
rect 476068 347244 476132 347308
rect 57100 347108 57164 347172
rect 60596 347108 60660 347172
rect 69796 347108 69860 347172
rect 192340 347108 192404 347172
rect 493364 347108 493428 347172
rect 460612 347032 460676 347036
rect 460612 346976 460626 347032
rect 460626 346976 460676 347032
rect 460612 346972 460676 346976
rect 465948 346972 466012 347036
rect 41828 346896 41892 346900
rect 41828 346840 41842 346896
rect 41842 346840 41892 346896
rect 41828 346836 41892 346840
rect 419580 346836 419644 346900
rect 54524 346700 54588 346764
rect 40540 346428 40604 346492
rect 18644 345204 18708 345268
rect 150940 335472 151004 335476
rect 150940 335416 150990 335472
rect 150990 335416 151004 335472
rect 150940 335412 151004 335416
rect 550956 335472 551020 335476
rect 550956 335416 551006 335472
rect 551006 335416 551020 335472
rect 550956 335412 551020 335416
rect 417740 278700 417804 278764
rect 417740 278156 417804 278220
rect 417556 260748 417620 260812
rect 417924 260748 417988 260812
rect 417556 259932 417620 259996
rect 191604 250412 191668 250476
rect 18828 249732 18892 249796
rect 93446 249792 93510 249796
rect 93446 249736 93490 249792
rect 93490 249736 93510 249792
rect 93446 249732 93510 249736
rect 95894 249792 95958 249796
rect 95894 249736 95938 249792
rect 95938 249736 95958 249792
rect 95894 249732 95958 249736
rect 98478 249732 98542 249796
rect 103510 249792 103574 249796
rect 103510 249736 103518 249792
rect 103518 249736 103574 249792
rect 103510 249732 103574 249736
rect 105958 249792 106022 249796
rect 105958 249736 106002 249792
rect 106002 249736 106022 249792
rect 105958 249732 106022 249736
rect 108542 249792 108606 249796
rect 108542 249736 108578 249792
rect 108578 249736 108606 249792
rect 108542 249732 108606 249736
rect 110990 249732 111054 249796
rect 468286 249732 468350 249796
rect 485966 249792 486030 249796
rect 485966 249736 486018 249792
rect 486018 249736 486030 249792
rect 485966 249732 486030 249736
rect 488278 249792 488342 249796
rect 488278 249736 488318 249792
rect 488318 249736 488342 249792
rect 488278 249732 488342 249736
rect 490998 249792 491062 249796
rect 490998 249736 491022 249792
rect 491022 249736 491062 249792
rect 490998 249732 491062 249736
rect 495894 249792 495958 249796
rect 495894 249736 495898 249792
rect 495898 249736 495954 249792
rect 495954 249736 495958 249792
rect 495894 249732 495958 249736
rect 498478 249792 498542 249796
rect 498478 249736 498530 249792
rect 498530 249736 498542 249792
rect 498478 249732 498542 249736
rect 500926 249792 500990 249796
rect 500926 249736 500958 249792
rect 500958 249736 500990 249792
rect 500926 249732 500990 249736
rect 503510 249792 503574 249796
rect 503510 249736 503534 249792
rect 503534 249736 503574 249792
rect 503510 249732 503574 249736
rect 50742 249656 50806 249660
rect 50742 249600 50802 249656
rect 50802 249600 50806 249656
rect 50742 249596 50806 249600
rect 53598 249656 53662 249660
rect 53598 249600 53654 249656
rect 53654 249600 53662 249656
rect 53598 249596 53662 249600
rect 56046 249656 56110 249660
rect 56046 249600 56102 249656
rect 56102 249600 56110 249656
rect 56046 249596 56110 249600
rect 58494 249656 58558 249660
rect 58494 249600 58530 249656
rect 58530 249600 58558 249656
rect 58494 249596 58558 249600
rect 113438 249656 113502 249660
rect 113438 249600 113454 249656
rect 113454 249600 113502 249656
rect 113438 249596 113502 249600
rect 115886 249656 115950 249660
rect 115886 249600 115902 249656
rect 115902 249600 115950 249656
rect 115886 249596 115950 249600
rect 120918 249656 120982 249660
rect 120918 249600 120962 249656
rect 120962 249600 120982 249656
rect 120918 249596 120982 249600
rect 461078 249596 461142 249660
rect 471006 249656 471070 249660
rect 471006 249600 471022 249656
rect 471022 249600 471070 249656
rect 471006 249596 471070 249600
rect 483518 249656 483582 249660
rect 483518 249600 483534 249656
rect 483534 249600 483582 249656
rect 483518 249596 483582 249600
rect 505958 249656 506022 249660
rect 505958 249600 505982 249656
rect 505982 249600 506022 249656
rect 505958 249596 506022 249600
rect 508542 249656 508606 249660
rect 508542 249600 508558 249656
rect 508558 249600 508606 249656
rect 508542 249596 508606 249600
rect 515886 249656 515950 249660
rect 515886 249600 515918 249656
rect 515918 249600 515950 249656
rect 515886 249596 515950 249600
rect 520918 249656 520982 249660
rect 520918 249600 520922 249656
rect 520922 249600 520978 249656
rect 520978 249600 520982 249656
rect 520918 249596 520982 249600
rect 418108 249460 418172 249524
rect 418844 249460 418908 249524
rect 476068 249460 476132 249524
rect 473676 249384 473740 249388
rect 473676 249328 473690 249384
rect 473690 249328 473740 249384
rect 473676 249324 473740 249328
rect 35940 248296 36004 248300
rect 35940 248240 35954 248296
rect 35954 248240 36004 248296
rect 35940 248236 36004 248240
rect 37044 248236 37108 248300
rect 39620 248236 39684 248300
rect 44220 248296 44284 248300
rect 44220 248240 44234 248296
rect 44234 248240 44284 248296
rect 44220 248236 44284 248240
rect 46612 248296 46676 248300
rect 46612 248240 46662 248296
rect 46662 248240 46676 248296
rect 46612 248236 46676 248240
rect 50108 248296 50172 248300
rect 50108 248240 50158 248296
rect 50158 248240 50172 248296
rect 50108 248236 50172 248240
rect 61148 248296 61212 248300
rect 61148 248240 61198 248296
rect 61198 248240 61212 248296
rect 61148 248236 61212 248240
rect 61700 248236 61764 248300
rect 62804 248236 62868 248300
rect 63540 248296 63604 248300
rect 63540 248240 63590 248296
rect 63590 248240 63604 248296
rect 63540 248236 63604 248240
rect 65196 248236 65260 248300
rect 65932 248296 65996 248300
rect 65932 248240 65982 248296
rect 65982 248240 65996 248296
rect 65932 248236 65996 248240
rect 68692 248236 68756 248300
rect 70900 248296 70964 248300
rect 70900 248240 70950 248296
rect 70950 248240 70964 248296
rect 70900 248236 70964 248240
rect 73660 248236 73724 248300
rect 78076 248236 78140 248300
rect 78444 248296 78508 248300
rect 78444 248240 78494 248296
rect 78494 248240 78508 248296
rect 78444 248236 78508 248240
rect 83596 248296 83660 248300
rect 83596 248240 83646 248296
rect 83646 248240 83660 248296
rect 83596 248236 83660 248240
rect 125916 248236 125980 248300
rect 443132 248296 443196 248300
rect 443132 248240 443182 248296
rect 443182 248240 443196 248296
rect 443132 248236 443196 248240
rect 448284 248236 448348 248300
rect 448652 248236 448716 248300
rect 450124 248296 450188 248300
rect 450124 248240 450174 248296
rect 450174 248240 450188 248296
rect 450124 248236 450188 248240
rect 450676 248236 450740 248300
rect 451228 248236 451292 248300
rect 453620 248236 453684 248300
rect 456196 248236 456260 248300
rect 462820 248236 462884 248300
rect 468708 248236 468772 248300
rect 38148 248100 38212 248164
rect 40540 248100 40604 248164
rect 41644 248100 41708 248164
rect 43116 248160 43180 248164
rect 43116 248104 43130 248160
rect 43130 248104 43180 248160
rect 43116 248100 43180 248104
rect 45324 248160 45388 248164
rect 45324 248104 45338 248160
rect 45338 248104 45388 248160
rect 45324 248100 45388 248104
rect 47532 248160 47596 248164
rect 47532 248104 47582 248160
rect 47582 248104 47596 248160
rect 47532 248100 47596 248104
rect 48452 248100 48516 248164
rect 478460 248100 478524 248164
rect 60596 247964 60660 248028
rect 48636 247888 48700 247892
rect 48636 247832 48686 247888
rect 48686 247832 48700 247888
rect 48636 247828 48700 247832
rect 58020 247888 58084 247892
rect 58020 247832 58070 247888
rect 58070 247832 58084 247888
rect 58020 247828 58084 247832
rect 59492 247888 59556 247892
rect 63908 247964 63972 248028
rect 79180 247964 79244 248028
rect 81020 248024 81084 248028
rect 81020 247968 81070 248024
rect 81070 247968 81084 248024
rect 81020 247964 81084 247968
rect 85988 248024 86052 248028
rect 85988 247968 86038 248024
rect 86038 247968 86052 248024
rect 85988 247964 86052 247968
rect 88196 248024 88260 248028
rect 88196 247968 88246 248024
rect 88246 247968 88260 248024
rect 88196 247964 88260 247968
rect 90956 248024 91020 248028
rect 90956 247968 91006 248024
rect 91006 247968 91020 248024
rect 90956 247964 91020 247968
rect 100892 247964 100956 248028
rect 118556 247964 118620 248028
rect 461716 247964 461780 248028
rect 465212 247964 465276 248028
rect 59492 247832 59506 247888
rect 59506 247832 59556 247888
rect 59492 247828 59556 247832
rect 66300 247888 66364 247892
rect 66300 247832 66314 247888
rect 66314 247832 66364 247888
rect 66300 247828 66364 247832
rect 67772 247888 67836 247892
rect 67772 247832 67786 247888
rect 67786 247832 67836 247888
rect 67772 247828 67836 247832
rect 68324 247888 68388 247892
rect 68324 247832 68374 247888
rect 68374 247832 68388 247888
rect 68324 247828 68388 247832
rect 76052 247888 76116 247892
rect 76052 247832 76102 247888
rect 76102 247832 76116 247888
rect 76052 247828 76116 247832
rect 123340 247828 123404 247892
rect 18828 247692 18892 247756
rect 75684 247692 75748 247756
rect 76972 247692 77036 247756
rect 458404 247692 458468 247756
rect 463556 247828 463620 247892
rect 463924 247828 463988 247892
rect 469812 247828 469876 247892
rect 474412 247828 474476 247892
rect 465948 247692 466012 247756
rect 467604 247692 467668 247756
rect 479196 247692 479260 247756
rect 18644 247556 18708 247620
rect 72188 247556 72252 247620
rect 455828 247616 455892 247620
rect 455828 247560 455878 247616
rect 455878 247560 455892 247616
rect 51396 247420 51460 247484
rect 69796 247420 69860 247484
rect 455828 247556 455892 247560
rect 460612 247556 460676 247620
rect 466316 247556 466380 247620
rect 471284 247556 471348 247620
rect 53420 247284 53484 247348
rect 71268 247284 71332 247348
rect 74396 247284 74460 247348
rect 437060 247284 437124 247348
rect 457116 247284 457180 247348
rect 475700 247420 475764 247484
rect 476988 247420 477052 247484
rect 459508 247344 459572 247348
rect 459508 247288 459522 247344
rect 459522 247288 459572 247344
rect 459508 247284 459572 247288
rect 472204 247284 472268 247348
rect 473308 247344 473372 247348
rect 473308 247288 473358 247344
rect 473358 247288 473372 247344
rect 473308 247284 473372 247288
rect 478092 247284 478156 247348
rect 73292 247148 73356 247212
rect 518388 247148 518452 247212
rect 52316 247072 52380 247076
rect 52316 247016 52366 247072
rect 52366 247016 52380 247072
rect 52316 247012 52380 247016
rect 54524 247012 54588 247076
rect 55812 247012 55876 247076
rect 57100 247012 57164 247076
rect 436140 247072 436204 247076
rect 436140 247016 436190 247072
rect 436190 247016 436204 247072
rect 436140 247012 436204 247016
rect 438164 247012 438228 247076
rect 439636 247012 439700 247076
rect 440556 247012 440620 247076
rect 441660 247072 441724 247076
rect 441660 247016 441674 247072
rect 441674 247016 441724 247072
rect 441660 247012 441724 247016
rect 444236 247072 444300 247076
rect 444236 247016 444286 247072
rect 444286 247016 444300 247072
rect 444236 247012 444300 247016
rect 445524 247012 445588 247076
rect 446628 247012 446692 247076
rect 447732 247012 447796 247076
rect 452332 247012 452396 247076
rect 453436 247012 453500 247076
rect 454540 247012 454604 247076
rect 458036 247072 458100 247076
rect 458036 247016 458086 247072
rect 458086 247016 458100 247072
rect 458036 247012 458100 247016
rect 480852 247012 480916 247076
rect 493364 247012 493428 247076
rect 511028 247012 511092 247076
rect 513420 247072 513484 247076
rect 513420 247016 513434 247072
rect 513434 247016 513484 247072
rect 513420 247012 513484 247016
rect 523356 247012 523420 247076
rect 525932 247012 525996 247076
rect 419948 238580 420012 238644
rect 419212 235860 419276 235924
rect 419580 235724 419644 235788
rect 550772 235104 550836 235108
rect 550772 235048 550822 235104
rect 550822 235048 550836 235104
rect 550772 235044 550836 235048
rect 150756 234636 150820 234700
rect 417924 179420 417988 179484
rect 417740 178196 417804 178260
rect 417556 159972 417620 160036
rect 19012 158068 19076 158132
rect 3372 149772 3436 149836
rect 458086 149832 458150 149836
rect 458086 149776 458142 149832
rect 458142 149776 458150 149832
rect 458086 149772 458150 149776
rect 478486 149832 478550 149836
rect 478486 149776 478510 149832
rect 478510 149776 478550 149832
rect 478486 149772 478550 149776
rect 480934 149832 480998 149836
rect 480934 149776 480958 149832
rect 480958 149776 480998 149832
rect 480934 149772 480998 149776
rect 483518 149832 483582 149836
rect 483518 149776 483534 149832
rect 483534 149776 483582 149832
rect 483518 149772 483582 149776
rect 485966 149832 486030 149836
rect 485966 149776 486018 149832
rect 486018 149776 486030 149832
rect 485966 149772 486030 149776
rect 440542 149636 440606 149700
rect 488278 149696 488342 149700
rect 488278 149640 488318 149696
rect 488318 149640 488342 149696
rect 488278 149636 488342 149640
rect 490998 149696 491062 149700
rect 490998 149640 491022 149696
rect 491022 149640 491062 149696
rect 490998 149636 491062 149640
rect 495894 149696 495958 149700
rect 495894 149640 495898 149696
rect 495898 149640 495954 149696
rect 495954 149640 495958 149696
rect 495894 149636 495958 149640
rect 503510 149696 503574 149700
rect 503510 149640 503534 149696
rect 503534 149640 503574 149696
rect 503510 149636 503574 149640
rect 48294 149560 48358 149564
rect 48294 149504 48318 149560
rect 48318 149504 48358 149560
rect 48294 149500 48358 149504
rect 50742 149560 50806 149564
rect 50742 149504 50802 149560
rect 50802 149504 50806 149560
rect 50742 149500 50806 149504
rect 56046 149560 56110 149564
rect 56046 149504 56102 149560
rect 56102 149504 56110 149560
rect 56046 149500 56110 149504
rect 58494 149560 58558 149564
rect 58494 149504 58530 149560
rect 58530 149504 58558 149560
rect 58494 149500 58558 149504
rect 60670 149560 60734 149564
rect 60670 149504 60702 149560
rect 60702 149504 60734 149560
rect 60670 149500 60734 149504
rect 71006 149500 71070 149564
rect 73590 149560 73654 149564
rect 73590 149504 73618 149560
rect 73618 149504 73654 149560
rect 73590 149500 73654 149504
rect 83518 149560 83582 149564
rect 83518 149504 83554 149560
rect 83554 149504 83582 149560
rect 83518 149500 83582 149504
rect 93446 149560 93510 149564
rect 93446 149504 93490 149560
rect 93490 149504 93510 149560
rect 93446 149500 93510 149504
rect 98478 149500 98542 149564
rect 103510 149560 103574 149564
rect 103510 149504 103518 149560
rect 103518 149504 103574 149560
rect 103510 149500 103574 149504
rect 113438 149560 113502 149564
rect 113438 149504 113454 149560
rect 113454 149504 113502 149560
rect 113438 149500 113502 149504
rect 115886 149560 115950 149564
rect 115886 149504 115902 149560
rect 115902 149504 115950 149560
rect 115886 149500 115950 149504
rect 120918 149560 120982 149564
rect 120918 149504 120962 149560
rect 120962 149504 120982 149560
rect 120918 149500 120982 149504
rect 441766 149500 441830 149564
rect 455910 149500 455974 149564
rect 461078 149500 461142 149564
rect 463526 149560 463590 149564
rect 463526 149504 463570 149560
rect 463570 149504 463590 149560
rect 463526 149500 463590 149504
rect 465974 149560 466038 149564
rect 465974 149504 465998 149560
rect 465998 149504 466038 149560
rect 465974 149500 466038 149504
rect 468286 149560 468350 149564
rect 468286 149504 468298 149560
rect 468298 149504 468350 149560
rect 468286 149500 468350 149504
rect 471006 149560 471070 149564
rect 471006 149504 471022 149560
rect 471022 149504 471070 149560
rect 471006 149500 471070 149504
rect 505958 149560 506022 149564
rect 505958 149504 505982 149560
rect 505982 149504 506022 149560
rect 505958 149500 506022 149504
rect 508542 149560 508606 149564
rect 508542 149504 508558 149560
rect 508558 149504 508606 149560
rect 508542 149500 508606 149504
rect 510990 149560 511054 149564
rect 510990 149504 511042 149560
rect 511042 149504 511054 149560
rect 510990 149500 511054 149504
rect 515886 149560 515950 149564
rect 515886 149504 515918 149560
rect 515918 149504 515950 149560
rect 515886 149500 515950 149504
rect 518470 149560 518534 149564
rect 518470 149504 518494 149560
rect 518494 149504 518534 149560
rect 518470 149500 518534 149504
rect 476068 149092 476132 149156
rect 53604 149016 53668 149020
rect 53604 148960 53654 149016
rect 53654 148960 53668 149016
rect 53604 148956 53668 148960
rect 76052 149016 76116 149020
rect 76052 148960 76102 149016
rect 76102 148960 76116 149016
rect 76052 148956 76116 148960
rect 85988 149016 86052 149020
rect 85988 148960 86038 149016
rect 86038 148960 86052 149016
rect 85988 148956 86052 148960
rect 123340 148956 123404 149020
rect 513420 149016 513484 149020
rect 513420 148960 513434 149016
rect 513434 148960 513484 149016
rect 513420 148956 513484 148960
rect 520964 149016 521028 149020
rect 520964 148960 520978 149016
rect 520978 148960 521028 149016
rect 520964 148956 521028 148960
rect 523356 149016 523420 149020
rect 523356 148960 523370 149016
rect 523370 148960 523420 149016
rect 523356 148956 523420 148960
rect 525932 149016 525996 149020
rect 525932 148960 525946 149016
rect 525946 148960 525996 149016
rect 525932 148956 525996 148960
rect 125916 148820 125980 148884
rect 459508 148744 459572 148748
rect 459508 148688 459522 148744
rect 459522 148688 459572 148744
rect 459508 148684 459572 148688
rect 419948 148276 420012 148340
rect 35940 147656 36004 147660
rect 35940 147600 35954 147656
rect 35954 147600 36004 147656
rect 35940 147596 36004 147600
rect 37044 147656 37108 147660
rect 37044 147600 37058 147656
rect 37058 147600 37108 147656
rect 37044 147596 37108 147600
rect 38148 147656 38212 147660
rect 38148 147600 38162 147656
rect 38162 147600 38212 147656
rect 38148 147596 38212 147600
rect 39620 147656 39684 147660
rect 39620 147600 39634 147656
rect 39634 147600 39684 147656
rect 39620 147596 39684 147600
rect 43116 147656 43180 147660
rect 43116 147600 43130 147656
rect 43130 147600 43180 147656
rect 43116 147596 43180 147600
rect 44220 147656 44284 147660
rect 44220 147600 44234 147656
rect 44234 147600 44284 147656
rect 44220 147596 44284 147600
rect 45324 147656 45388 147660
rect 45324 147600 45338 147656
rect 45338 147600 45388 147656
rect 45324 147596 45388 147600
rect 46612 147656 46676 147660
rect 46612 147600 46626 147656
rect 46626 147600 46676 147656
rect 46612 147596 46676 147600
rect 47716 147656 47780 147660
rect 47716 147600 47730 147656
rect 47730 147600 47780 147656
rect 47716 147596 47780 147600
rect 48636 147656 48700 147660
rect 48636 147600 48686 147656
rect 48686 147600 48700 147656
rect 48636 147596 48700 147600
rect 50108 147656 50172 147660
rect 50108 147600 50158 147656
rect 50158 147600 50172 147656
rect 50108 147596 50172 147600
rect 51396 147656 51460 147660
rect 51396 147600 51446 147656
rect 51446 147600 51460 147656
rect 51396 147596 51460 147600
rect 52316 147656 52380 147660
rect 52316 147600 52330 147656
rect 52330 147600 52380 147656
rect 52316 147596 52380 147600
rect 53420 147656 53484 147660
rect 53420 147600 53434 147656
rect 53434 147600 53484 147656
rect 53420 147596 53484 147600
rect 54524 147596 54588 147660
rect 55996 147656 56060 147660
rect 55996 147600 56046 147656
rect 56046 147600 56060 147656
rect 55996 147596 56060 147600
rect 58020 147656 58084 147660
rect 58020 147600 58070 147656
rect 58070 147600 58084 147656
rect 58020 147596 58084 147600
rect 59492 147656 59556 147660
rect 59492 147600 59542 147656
rect 59542 147600 59556 147656
rect 59492 147596 59556 147600
rect 61700 147656 61764 147660
rect 61700 147600 61714 147656
rect 61714 147600 61764 147656
rect 61700 147596 61764 147600
rect 62804 147656 62868 147660
rect 62804 147600 62818 147656
rect 62818 147600 62868 147656
rect 62804 147596 62868 147600
rect 63540 147656 63604 147660
rect 63540 147600 63590 147656
rect 63590 147600 63604 147656
rect 63540 147596 63604 147600
rect 63908 147656 63972 147660
rect 63908 147600 63922 147656
rect 63922 147600 63972 147656
rect 63908 147596 63972 147600
rect 65196 147656 65260 147660
rect 65196 147600 65210 147656
rect 65210 147600 65260 147656
rect 65196 147596 65260 147600
rect 66116 147656 66180 147660
rect 66116 147600 66166 147656
rect 66166 147600 66180 147656
rect 66116 147596 66180 147600
rect 66300 147656 66364 147660
rect 66300 147600 66350 147656
rect 66350 147600 66364 147656
rect 66300 147596 66364 147600
rect 67588 147656 67652 147660
rect 67588 147600 67638 147656
rect 67638 147600 67652 147656
rect 67588 147596 67652 147600
rect 68140 147596 68204 147660
rect 68692 147596 68756 147660
rect 69796 147656 69860 147660
rect 69796 147600 69810 147656
rect 69810 147600 69860 147656
rect 69796 147596 69860 147600
rect 72188 147656 72252 147660
rect 72188 147600 72202 147656
rect 72202 147600 72252 147656
rect 72188 147596 72252 147600
rect 73292 147656 73356 147660
rect 73292 147600 73306 147656
rect 73306 147600 73356 147656
rect 73292 147596 73356 147600
rect 74396 147596 74460 147660
rect 75684 147656 75748 147660
rect 75684 147600 75698 147656
rect 75698 147600 75748 147656
rect 75684 147596 75748 147600
rect 76972 147656 77036 147660
rect 76972 147600 76986 147656
rect 76986 147600 77036 147656
rect 76972 147596 77036 147600
rect 78076 147656 78140 147660
rect 78076 147600 78090 147656
rect 78090 147600 78140 147656
rect 78076 147596 78140 147600
rect 78444 147656 78508 147660
rect 78444 147600 78494 147656
rect 78494 147600 78508 147656
rect 78444 147596 78508 147600
rect 79180 147656 79244 147660
rect 79180 147600 79194 147656
rect 79194 147600 79244 147656
rect 79180 147596 79244 147600
rect 81020 147656 81084 147660
rect 81020 147600 81070 147656
rect 81070 147600 81084 147656
rect 81020 147596 81084 147600
rect 88196 147656 88260 147660
rect 88196 147600 88246 147656
rect 88246 147600 88260 147656
rect 88196 147596 88260 147600
rect 90956 147656 91020 147660
rect 90956 147600 91006 147656
rect 91006 147600 91020 147656
rect 90956 147596 91020 147600
rect 95924 147656 95988 147660
rect 95924 147600 95974 147656
rect 95974 147600 95988 147656
rect 95924 147596 95988 147600
rect 100892 147656 100956 147660
rect 100892 147600 100942 147656
rect 100942 147600 100956 147656
rect 100892 147596 100956 147600
rect 106044 147656 106108 147660
rect 106044 147600 106094 147656
rect 106094 147600 106108 147656
rect 106044 147596 106108 147600
rect 108620 147596 108684 147660
rect 111012 147596 111076 147660
rect 436140 147656 436204 147660
rect 436140 147600 436154 147656
rect 436154 147600 436204 147656
rect 436140 147596 436204 147600
rect 437060 147656 437124 147660
rect 437060 147600 437074 147656
rect 437074 147600 437124 147656
rect 437060 147596 437124 147600
rect 437980 147656 438044 147660
rect 437980 147600 437994 147656
rect 437994 147600 438044 147656
rect 437980 147596 438044 147600
rect 439636 147656 439700 147660
rect 439636 147600 439650 147656
rect 439650 147600 439700 147656
rect 439636 147596 439700 147600
rect 443132 147656 443196 147660
rect 443132 147600 443146 147656
rect 443146 147600 443196 147656
rect 443132 147596 443196 147600
rect 444236 147656 444300 147660
rect 444236 147600 444250 147656
rect 444250 147600 444300 147656
rect 444236 147596 444300 147600
rect 445340 147656 445404 147660
rect 445340 147600 445354 147656
rect 445354 147600 445404 147656
rect 445340 147596 445404 147600
rect 446444 147656 446508 147660
rect 446444 147600 446458 147656
rect 446458 147600 446508 147656
rect 446444 147596 446508 147600
rect 447364 147596 447428 147660
rect 448284 147656 448348 147660
rect 448284 147600 448298 147656
rect 448298 147600 448348 147656
rect 448284 147596 448348 147600
rect 448652 147596 448716 147660
rect 450124 147596 450188 147660
rect 450676 147656 450740 147660
rect 450676 147600 450690 147656
rect 450690 147600 450740 147656
rect 450676 147596 450740 147600
rect 451228 147656 451292 147660
rect 451228 147600 451278 147656
rect 451278 147600 451292 147656
rect 451228 147596 451292 147600
rect 452332 147596 452396 147660
rect 453436 147656 453500 147660
rect 453436 147600 453450 147656
rect 453450 147600 453500 147656
rect 453436 147596 453500 147600
rect 453620 147656 453684 147660
rect 453620 147600 453634 147656
rect 453634 147600 453684 147656
rect 453620 147596 453684 147600
rect 454540 147656 454604 147660
rect 454540 147600 454590 147656
rect 454590 147600 454604 147656
rect 454540 147596 454604 147600
rect 456012 147656 456076 147660
rect 456012 147600 456026 147656
rect 456026 147600 456076 147656
rect 456012 147596 456076 147600
rect 458404 147656 458468 147660
rect 458404 147600 458418 147656
rect 458418 147600 458468 147656
rect 458404 147596 458468 147600
rect 461716 147656 461780 147660
rect 461716 147600 461730 147656
rect 461730 147600 461780 147656
rect 461716 147596 461780 147600
rect 462820 147656 462884 147660
rect 462820 147600 462834 147656
rect 462834 147600 462884 147656
rect 462820 147596 462884 147600
rect 463924 147656 463988 147660
rect 463924 147600 463938 147656
rect 463938 147600 463988 147656
rect 463924 147596 463988 147600
rect 465212 147656 465276 147660
rect 465212 147600 465226 147656
rect 465226 147600 465276 147656
rect 465212 147596 465276 147600
rect 466316 147656 466380 147660
rect 466316 147600 466330 147656
rect 466330 147600 466380 147656
rect 466316 147596 466380 147600
rect 467604 147656 467668 147660
rect 467604 147600 467618 147656
rect 467618 147600 467668 147656
rect 467604 147596 467668 147600
rect 468708 147656 468772 147660
rect 468708 147600 468722 147656
rect 468722 147600 468772 147656
rect 468708 147596 468772 147600
rect 469812 147656 469876 147660
rect 469812 147600 469826 147656
rect 469826 147600 469876 147656
rect 469812 147596 469876 147600
rect 471100 147656 471164 147660
rect 471100 147600 471114 147656
rect 471114 147600 471164 147656
rect 471100 147596 471164 147600
rect 472204 147656 472268 147660
rect 472204 147600 472218 147656
rect 472218 147600 472268 147656
rect 472204 147596 472268 147600
rect 473308 147656 473372 147660
rect 473308 147600 473358 147656
rect 473358 147600 473372 147656
rect 473308 147596 473372 147600
rect 474412 147596 474476 147660
rect 476988 147656 477052 147660
rect 476988 147600 477002 147656
rect 477002 147600 477052 147656
rect 476988 147596 477052 147600
rect 478092 147656 478156 147660
rect 478092 147600 478106 147656
rect 478106 147600 478156 147656
rect 478092 147596 478156 147600
rect 18644 147460 18708 147524
rect 41828 147460 41892 147524
rect 118556 147460 118620 147524
rect 500908 147460 500972 147524
rect 40540 147324 40604 147388
rect 61148 147324 61212 147388
rect 493364 147324 493428 147388
rect 56916 147188 56980 147252
rect 71084 147248 71148 147252
rect 71084 147192 71098 147248
rect 71098 147192 71148 147248
rect 71084 147188 71148 147192
rect 419396 147188 419460 147252
rect 473492 147188 473556 147252
rect 456932 147052 456996 147116
rect 460612 146916 460676 146980
rect 479196 147052 479260 147116
rect 18828 146840 18892 146844
rect 18828 146784 18842 146840
rect 18842 146784 18892 146840
rect 18828 146780 18892 146784
rect 419212 146780 419276 146844
rect 456932 146780 456996 146844
rect 475516 146780 475580 146844
rect 498516 146508 498580 146572
rect 551508 136444 551572 136508
rect 151124 135764 151188 135828
rect 417924 79868 417988 79932
rect 417740 78100 417804 78164
rect 417556 59876 417620 59940
rect 19196 57972 19260 58036
rect 53462 49872 53526 49876
rect 53462 49816 53470 49872
rect 53470 49816 53526 49872
rect 53462 49812 53526 49816
rect 60670 49872 60734 49876
rect 60670 49816 60702 49872
rect 60702 49816 60734 49872
rect 60670 49812 60734 49816
rect 456998 49872 457062 49876
rect 456998 49816 457038 49872
rect 457038 49816 457062 49872
rect 456998 49812 457062 49816
rect 458086 49872 458150 49876
rect 458086 49816 458142 49872
rect 458142 49816 458150 49872
rect 458086 49812 458150 49816
rect 478486 49872 478550 49876
rect 478486 49816 478510 49872
rect 478510 49816 478550 49872
rect 478486 49812 478550 49816
rect 480934 49872 480998 49876
rect 480934 49816 480958 49872
rect 480958 49816 480998 49872
rect 480934 49812 480998 49816
rect 90998 49736 91062 49740
rect 90998 49680 91006 49736
rect 91006 49680 91062 49736
rect 90998 49676 91062 49680
rect 95894 49736 95958 49740
rect 95894 49680 95938 49736
rect 95938 49680 95958 49736
rect 95894 49676 95958 49680
rect 473318 49736 473382 49740
rect 473318 49680 473358 49736
rect 473358 49680 473382 49736
rect 473318 49676 473382 49680
rect 488278 49736 488342 49740
rect 488278 49680 488318 49736
rect 488318 49680 488342 49736
rect 488278 49676 488342 49680
rect 495894 49736 495958 49740
rect 495894 49680 495898 49736
rect 495898 49680 495954 49736
rect 495954 49680 495958 49736
rect 495894 49676 495958 49680
rect 503510 49736 503574 49740
rect 503510 49680 503534 49736
rect 503534 49680 503574 49736
rect 503510 49676 503574 49680
rect 48294 49600 48358 49604
rect 48294 49544 48318 49600
rect 48318 49544 48358 49600
rect 48294 49540 48358 49544
rect 50742 49600 50806 49604
rect 50742 49544 50802 49600
rect 50802 49544 50806 49600
rect 50742 49540 50806 49544
rect 53598 49600 53662 49604
rect 53598 49544 53654 49600
rect 53654 49544 53662 49600
rect 53598 49540 53662 49544
rect 56046 49600 56110 49604
rect 56046 49544 56102 49600
rect 56102 49544 56110 49600
rect 56046 49540 56110 49544
rect 58494 49600 58558 49604
rect 58494 49544 58530 49600
rect 58530 49544 58558 49600
rect 58494 49540 58558 49544
rect 80934 49600 80998 49604
rect 80934 49544 80978 49600
rect 80978 49544 80998 49600
rect 80934 49540 80998 49544
rect 83518 49600 83582 49604
rect 83518 49544 83554 49600
rect 83554 49544 83582 49600
rect 83518 49540 83582 49544
rect 85966 49540 86030 49604
rect 88278 49600 88342 49604
rect 88278 49544 88302 49600
rect 88302 49544 88342 49600
rect 88278 49540 88342 49544
rect 98478 49540 98542 49604
rect 103510 49600 103574 49604
rect 103510 49544 103518 49600
rect 103518 49544 103574 49600
rect 103510 49540 103574 49544
rect 105958 49600 106022 49604
rect 105958 49544 106002 49600
rect 106002 49544 106022 49600
rect 105958 49540 106022 49544
rect 120918 49540 120982 49604
rect 490998 49540 491062 49604
rect 493446 49600 493510 49604
rect 493446 49544 493470 49600
rect 493470 49544 493510 49600
rect 493446 49540 493510 49544
rect 498478 49600 498542 49604
rect 498478 49544 498530 49600
rect 498530 49544 498542 49600
rect 498478 49540 498542 49544
rect 500926 49600 500990 49604
rect 500926 49544 500958 49600
rect 500958 49544 500990 49600
rect 500926 49540 500990 49544
rect 505958 49600 506022 49604
rect 505958 49544 505982 49600
rect 505982 49544 506022 49600
rect 505958 49540 506022 49544
rect 508542 49600 508606 49604
rect 508542 49544 508558 49600
rect 508558 49544 508606 49600
rect 508542 49540 508606 49544
rect 510990 49600 511054 49604
rect 510990 49544 511042 49600
rect 511042 49544 511054 49600
rect 510990 49540 511054 49544
rect 513438 49540 513502 49604
rect 515886 49600 515950 49604
rect 515886 49544 515918 49600
rect 515918 49544 515950 49600
rect 515886 49540 515950 49544
rect 520918 49600 520982 49604
rect 520918 49544 520922 49600
rect 520922 49544 520978 49600
rect 520978 49544 520982 49600
rect 520918 49540 520982 49544
rect 525950 49540 526014 49604
rect 113404 49404 113468 49468
rect 486004 49404 486068 49468
rect 483428 49268 483492 49332
rect 418660 49132 418724 49196
rect 460980 49132 461044 49196
rect 419948 48996 420012 49060
rect 459508 49056 459572 49060
rect 459508 49000 459522 49056
rect 459522 49000 459572 49056
rect 459508 48996 459572 49000
rect 37044 48180 37108 48244
rect 43116 48240 43180 48244
rect 43116 48184 43166 48240
rect 43166 48184 43180 48240
rect 43116 48180 43180 48184
rect 44220 48240 44284 48244
rect 44220 48184 44234 48240
rect 44234 48184 44284 48240
rect 44220 48180 44284 48184
rect 45324 48240 45388 48244
rect 45324 48184 45374 48240
rect 45374 48184 45388 48240
rect 45324 48180 45388 48184
rect 46612 48240 46676 48244
rect 46612 48184 46626 48240
rect 46626 48184 46676 48240
rect 46612 48180 46676 48184
rect 47532 48240 47596 48244
rect 47532 48184 47582 48240
rect 47582 48184 47596 48240
rect 47532 48180 47596 48184
rect 48636 48240 48700 48244
rect 48636 48184 48686 48240
rect 48686 48184 48700 48240
rect 48636 48180 48700 48184
rect 50108 48180 50172 48244
rect 51396 48240 51460 48244
rect 51396 48184 51446 48240
rect 51446 48184 51460 48240
rect 51396 48180 51460 48184
rect 52316 48240 52380 48244
rect 52316 48184 52366 48240
rect 52366 48184 52380 48240
rect 52316 48180 52380 48184
rect 54524 48240 54588 48244
rect 54524 48184 54574 48240
rect 54574 48184 54588 48240
rect 54524 48180 54588 48184
rect 55812 48240 55876 48244
rect 55812 48184 55862 48240
rect 55862 48184 55876 48240
rect 55812 48180 55876 48184
rect 58020 48240 58084 48244
rect 58020 48184 58034 48240
rect 58034 48184 58084 48240
rect 58020 48180 58084 48184
rect 59492 48240 59556 48244
rect 59492 48184 59542 48240
rect 59542 48184 59556 48240
rect 59492 48180 59556 48184
rect 61148 48240 61212 48244
rect 61148 48184 61198 48240
rect 61198 48184 61212 48240
rect 61148 48180 61212 48184
rect 61700 48180 61764 48244
rect 62804 48180 62868 48244
rect 63540 48180 63604 48244
rect 65196 48180 65260 48244
rect 65932 48240 65996 48244
rect 65932 48184 65982 48240
rect 65982 48184 65996 48240
rect 65932 48180 65996 48184
rect 66300 48240 66364 48244
rect 66300 48184 66314 48240
rect 66314 48184 66364 48240
rect 66300 48180 66364 48184
rect 67588 48240 67652 48244
rect 67588 48184 67638 48240
rect 67638 48184 67652 48240
rect 67588 48180 67652 48184
rect 68324 48240 68388 48244
rect 68324 48184 68374 48240
rect 68374 48184 68388 48240
rect 68324 48180 68388 48184
rect 68692 48180 68756 48244
rect 69796 48240 69860 48244
rect 69796 48184 69810 48240
rect 69810 48184 69860 48240
rect 69796 48180 69860 48184
rect 70900 48180 70964 48244
rect 72188 48180 72252 48244
rect 73292 48240 73356 48244
rect 73292 48184 73306 48240
rect 73306 48184 73356 48240
rect 73292 48180 73356 48184
rect 73660 48180 73724 48244
rect 74396 48240 74460 48244
rect 74396 48184 74410 48240
rect 74410 48184 74460 48240
rect 74396 48180 74460 48184
rect 76052 48240 76116 48244
rect 76052 48184 76102 48240
rect 76102 48184 76116 48240
rect 76052 48180 76116 48184
rect 76972 48180 77036 48244
rect 78076 48240 78140 48244
rect 78076 48184 78090 48240
rect 78090 48184 78140 48240
rect 78076 48180 78140 48184
rect 78444 48240 78508 48244
rect 78444 48184 78494 48240
rect 78494 48184 78508 48240
rect 78444 48180 78508 48184
rect 93532 48240 93596 48244
rect 93532 48184 93582 48240
rect 93582 48184 93596 48240
rect 93532 48180 93596 48184
rect 100892 48240 100956 48244
rect 100892 48184 100942 48240
rect 100942 48184 100956 48240
rect 100892 48180 100956 48184
rect 108620 48180 108684 48244
rect 111012 48180 111076 48244
rect 115796 48240 115860 48244
rect 115796 48184 115846 48240
rect 115846 48184 115860 48240
rect 115796 48180 115860 48184
rect 118556 48240 118620 48244
rect 118556 48184 118606 48240
rect 118606 48184 118620 48240
rect 118556 48180 118620 48184
rect 125916 48240 125980 48244
rect 125916 48184 125966 48240
rect 125966 48184 125980 48240
rect 125916 48180 125980 48184
rect 436140 48240 436204 48244
rect 436140 48184 436154 48240
rect 436154 48184 436204 48240
rect 436140 48180 436204 48184
rect 437060 48240 437124 48244
rect 437060 48184 437074 48240
rect 437074 48184 437124 48240
rect 437060 48180 437124 48184
rect 438164 48240 438228 48244
rect 438164 48184 438178 48240
rect 438178 48184 438228 48240
rect 438164 48180 438228 48184
rect 439636 48240 439700 48244
rect 439636 48184 439650 48240
rect 439650 48184 439700 48240
rect 439636 48180 439700 48184
rect 443132 48240 443196 48244
rect 443132 48184 443146 48240
rect 443146 48184 443196 48240
rect 443132 48180 443196 48184
rect 444236 48240 444300 48244
rect 444236 48184 444286 48240
rect 444286 48184 444300 48240
rect 444236 48180 444300 48184
rect 448284 48240 448348 48244
rect 448284 48184 448298 48240
rect 448298 48184 448348 48240
rect 448284 48180 448348 48184
rect 450676 48240 450740 48244
rect 450676 48184 450690 48240
rect 450690 48184 450740 48240
rect 450676 48180 450740 48184
rect 453620 48240 453684 48244
rect 453620 48184 453634 48240
rect 453634 48184 453684 48240
rect 453620 48180 453684 48184
rect 454540 48240 454604 48244
rect 454540 48184 454590 48240
rect 454590 48184 454604 48240
rect 454540 48180 454604 48184
rect 455644 48180 455708 48244
rect 458404 48240 458468 48244
rect 458404 48184 458418 48240
rect 458418 48184 458468 48240
rect 458404 48180 458468 48184
rect 461716 48240 461780 48244
rect 461716 48184 461730 48240
rect 461730 48184 461780 48240
rect 461716 48180 461780 48184
rect 462820 48240 462884 48244
rect 462820 48184 462834 48240
rect 462834 48184 462884 48240
rect 462820 48180 462884 48184
rect 463556 48240 463620 48244
rect 463556 48184 463570 48240
rect 463570 48184 463620 48240
rect 463556 48180 463620 48184
rect 463924 48240 463988 48244
rect 463924 48184 463938 48240
rect 463938 48184 463988 48240
rect 463924 48180 463988 48184
rect 465212 48240 465276 48244
rect 465212 48184 465226 48240
rect 465226 48184 465276 48240
rect 465212 48180 465276 48184
rect 465948 48240 466012 48244
rect 465948 48184 465962 48240
rect 465962 48184 466012 48240
rect 465948 48180 466012 48184
rect 466316 48240 466380 48244
rect 466316 48184 466330 48240
rect 466330 48184 466380 48240
rect 466316 48180 466380 48184
rect 467604 48240 467668 48244
rect 467604 48184 467618 48240
rect 467618 48184 467668 48240
rect 467604 48180 467668 48184
rect 468340 48240 468404 48244
rect 468340 48184 468354 48240
rect 468354 48184 468404 48240
rect 468340 48180 468404 48184
rect 468708 48240 468772 48244
rect 468708 48184 468722 48240
rect 468722 48184 468772 48240
rect 468708 48180 468772 48184
rect 469812 48180 469876 48244
rect 470916 48240 470980 48244
rect 470916 48184 470930 48240
rect 470930 48184 470980 48240
rect 470916 48180 470980 48184
rect 471284 48240 471348 48244
rect 471284 48184 471298 48240
rect 471298 48184 471348 48240
rect 471284 48180 471348 48184
rect 472204 48240 472268 48244
rect 472204 48184 472218 48240
rect 472218 48184 472268 48240
rect 472204 48180 472268 48184
rect 474412 48240 474476 48244
rect 474412 48184 474426 48240
rect 474426 48184 474476 48240
rect 474412 48180 474476 48184
rect 475700 48240 475764 48244
rect 475700 48184 475714 48240
rect 475714 48184 475764 48240
rect 475700 48180 475764 48184
rect 476988 48240 477052 48244
rect 476988 48184 477002 48240
rect 477002 48184 477052 48240
rect 476988 48180 477052 48184
rect 478092 48240 478156 48244
rect 478092 48184 478106 48240
rect 478106 48184 478156 48240
rect 478092 48180 478156 48184
rect 40540 48044 40604 48108
rect 41828 48044 41892 48108
rect 63908 48104 63972 48108
rect 63908 48048 63922 48104
rect 63922 48048 63972 48104
rect 63908 48044 63972 48048
rect 71084 48104 71148 48108
rect 71084 48048 71098 48104
rect 71098 48048 71148 48104
rect 71084 48044 71148 48048
rect 123340 48044 123404 48108
rect 389220 48044 389284 48108
rect 419396 48044 419460 48108
rect 440556 48044 440620 48108
rect 445340 48104 445404 48108
rect 445340 48048 445354 48104
rect 445354 48048 445404 48104
rect 445340 48044 445404 48048
rect 446444 48104 446508 48108
rect 446444 48048 446458 48104
rect 446458 48048 446508 48104
rect 446444 48044 446508 48048
rect 448652 48044 448716 48108
rect 39620 47908 39684 47972
rect 38516 47772 38580 47836
rect 18644 47636 18708 47700
rect 452332 48104 452396 48108
rect 452332 48048 452346 48104
rect 452346 48048 452396 48104
rect 452332 48044 452396 48048
rect 453436 48044 453500 48108
rect 79180 47908 79244 47972
rect 475884 47908 475948 47972
rect 473308 47772 473372 47836
rect 415900 47636 415964 47700
rect 455828 47636 455892 47700
rect 460612 47636 460676 47700
rect 479196 47636 479260 47700
rect 35940 47500 36004 47564
rect 57100 47560 57164 47564
rect 57100 47504 57114 47560
rect 57114 47504 57164 47560
rect 57100 47500 57164 47504
rect 75684 47500 75748 47564
rect 419212 47500 419276 47564
rect 447548 47560 447612 47564
rect 447548 47504 447562 47560
rect 447562 47504 447612 47560
rect 447548 47500 447612 47504
rect 442028 47364 442092 47428
rect 450124 47424 450188 47428
rect 450124 47368 450138 47424
rect 450138 47368 450188 47424
rect 450124 47364 450188 47368
rect 451228 47424 451292 47428
rect 451228 47368 451278 47424
rect 451278 47368 451292 47424
rect 451228 47364 451292 47368
rect 523356 47228 523420 47292
rect 518388 47092 518452 47156
rect 193812 31724 193876 31788
rect 193996 19348 194060 19412
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 3371 466580 3437 466581
rect 3371 466516 3372 466580
rect 3436 466516 3437 466580
rect 3371 466515 3437 466516
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 3374 149837 3434 466515
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 3371 149836 3437 149837
rect 3371 149772 3372 149836
rect 3436 149772 3437 149836
rect 3371 149771 3437 149772
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 19195 455700 19261 455701
rect 19195 455636 19196 455700
rect 19260 455636 19261 455700
rect 19195 455635 19261 455636
rect 19011 453388 19077 453389
rect 19011 453324 19012 453388
rect 19076 453324 19077 453388
rect 19011 453323 19077 453324
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 18643 345268 18709 345269
rect 18643 345204 18644 345268
rect 18708 345204 18709 345268
rect 18643 345203 18709 345204
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 18646 247621 18706 345203
rect 18827 249796 18893 249797
rect 18827 249732 18828 249796
rect 18892 249732 18893 249796
rect 18827 249731 18893 249732
rect 18830 247757 18890 249731
rect 18827 247756 18893 247757
rect 18827 247692 18828 247756
rect 18892 247692 18893 247756
rect 18827 247691 18893 247692
rect 18643 247620 18709 247621
rect 18643 247556 18644 247620
rect 18708 247556 18709 247620
rect 18643 247555 18709 247556
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 18646 147525 18706 247555
rect 18643 147524 18709 147525
rect 18643 147460 18644 147524
rect 18708 147460 18709 147524
rect 18643 147459 18709 147460
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 18646 47701 18706 147459
rect 18830 146845 18890 247691
rect 19014 158133 19074 453323
rect 19011 158132 19077 158133
rect 19011 158068 19012 158132
rect 19076 158068 19077 158132
rect 19011 158067 19077 158068
rect 18827 146844 18893 146845
rect 18827 146780 18828 146844
rect 18892 146780 18893 146844
rect 18827 146779 18893 146780
rect 19198 58037 19258 455635
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 435244 21014 453498
rect 24114 493774 24734 500068
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 435244 24734 457218
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 435244 28454 460938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435244 38414 470898
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 435244 42134 438618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 435244 45854 442338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 435244 49574 446058
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52674 558334 53294 593778
rect 56394 598054 57014 633498
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52674 522334 53294 557778
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52674 486334 53294 521778
rect 56394 526054 57014 561498
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52674 435244 53294 449778
rect 56394 490054 57014 525498
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 435244 57014 453498
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 678961 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 678961 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 678961 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 678961 85574 698058
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 678961 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 678961 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 678961 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 678961 121574 698058
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 678961 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 678961 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 601774 60734 637218
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 60114 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 60734 601774
rect 60114 601454 60734 601538
rect 60114 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 60734 601454
rect 60114 565774 60734 601218
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 60114 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 60734 565774
rect 60114 565454 60734 565538
rect 60114 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 60734 565454
rect 60114 529774 60734 565218
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 60114 493774 60734 529218
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 60114 435244 60734 457218
rect 63834 497494 64454 501375
rect 63834 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 64454 497494
rect 63834 497174 64454 497258
rect 63834 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 64454 497174
rect 63834 461494 64454 496938
rect 63834 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 64454 461494
rect 63834 461174 64454 461258
rect 63834 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 64454 461174
rect 63834 435244 64454 460938
rect 73794 471454 74414 501375
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435244 74414 470898
rect 77514 475174 78134 501375
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 435244 78134 438618
rect 81234 478894 81854 501375
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 435244 81854 442338
rect 84954 482614 85574 501375
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 435244 85574 446058
rect 88674 486334 89294 501375
rect 88674 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 89294 486334
rect 88674 486014 89294 486098
rect 88674 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 89294 486014
rect 88674 450334 89294 485778
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 88674 435244 89294 449778
rect 92394 490054 93014 501375
rect 92394 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 93014 490054
rect 92394 489734 93014 489818
rect 92394 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 93014 489734
rect 92394 454054 93014 489498
rect 92394 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 93014 454054
rect 92394 453734 93014 453818
rect 92394 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 93014 453734
rect 92394 435244 93014 453498
rect 96114 493774 96734 501375
rect 96114 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 96734 493774
rect 96114 493454 96734 493538
rect 96114 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 96734 493454
rect 96114 457774 96734 493218
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 96114 435244 96734 457218
rect 99834 497494 100454 501375
rect 99834 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 100454 497494
rect 99834 497174 100454 497258
rect 99834 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 100454 497174
rect 99834 461494 100454 496938
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 99834 435244 100454 460938
rect 109794 471454 110414 501375
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435244 110414 470898
rect 113514 475174 114134 501375
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 435244 114134 438618
rect 117234 478894 117854 501375
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 435244 117854 442338
rect 120954 482614 121574 501375
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 435244 121574 446058
rect 124674 486334 125294 501375
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 124674 450334 125294 485778
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 435244 125294 449778
rect 128394 490054 129014 501375
rect 128394 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 129014 490054
rect 128394 489734 129014 489818
rect 128394 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 129014 489734
rect 128394 454054 129014 489498
rect 128394 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 129014 454054
rect 128394 453734 129014 453818
rect 128394 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 129014 453734
rect 128394 435244 129014 453498
rect 132114 493774 132734 501375
rect 132114 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 132734 493774
rect 132114 493454 132734 493538
rect 132114 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 132734 493454
rect 132114 457774 132734 493218
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 132114 435244 132734 457218
rect 135834 497494 136454 501375
rect 135834 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 136454 497494
rect 135834 497174 136454 497258
rect 135834 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 136454 497174
rect 135834 461494 136454 496938
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 135834 435244 136454 460938
rect 145794 471454 146414 501375
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435244 146414 470898
rect 149514 475174 150134 501375
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 435244 150134 438618
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 150939 435300 151005 435301
rect 150939 435236 150940 435300
rect 151004 435236 151005 435300
rect 153234 435244 153854 442338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 435244 157574 446058
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 160674 594334 161294 629778
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 160674 558334 161294 593778
rect 164394 598054 165014 633498
rect 164394 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 165014 598054
rect 164394 597734 165014 597818
rect 164394 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 165014 597734
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 160674 522334 161294 557778
rect 164394 562054 165014 597498
rect 164394 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 165014 562054
rect 164394 561734 165014 561818
rect 164394 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 165014 561734
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 160674 486334 161294 521778
rect 164394 526054 165014 561498
rect 164394 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 165014 526054
rect 164394 525734 165014 525818
rect 164394 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 165014 525734
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 160674 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 161294 486334
rect 160674 486014 161294 486098
rect 160674 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 161294 486014
rect 160674 450334 161294 485778
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 150939 435235 151005 435236
rect 150942 433530 151002 435235
rect 150840 433470 151002 433530
rect 150840 433202 150900 433470
rect 160674 414334 161294 449778
rect 160674 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 161294 414334
rect 160674 414014 161294 414098
rect 160674 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 161294 414014
rect 20272 403174 20620 403206
rect 20272 402938 20328 403174
rect 20564 402938 20620 403174
rect 20272 402854 20620 402938
rect 20272 402618 20328 402854
rect 20564 402618 20620 402854
rect 20272 402586 20620 402618
rect 156000 403174 156348 403206
rect 156000 402938 156056 403174
rect 156292 402938 156348 403174
rect 156000 402854 156348 402938
rect 156000 402618 156056 402854
rect 156292 402618 156348 402854
rect 156000 402586 156348 402618
rect 20952 399454 21300 399486
rect 20952 399218 21008 399454
rect 21244 399218 21300 399454
rect 20952 399134 21300 399218
rect 20952 398898 21008 399134
rect 21244 398898 21300 399134
rect 20952 398866 21300 398898
rect 155320 399454 155668 399486
rect 155320 399218 155376 399454
rect 155612 399218 155668 399454
rect 155320 399134 155668 399218
rect 155320 398898 155376 399134
rect 155612 398898 155668 399134
rect 155320 398866 155668 398898
rect 160674 378334 161294 413778
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 20272 367174 20620 367206
rect 20272 366938 20328 367174
rect 20564 366938 20620 367174
rect 20272 366854 20620 366938
rect 20272 366618 20328 366854
rect 20564 366618 20620 366854
rect 20272 366586 20620 366618
rect 156000 367174 156348 367206
rect 156000 366938 156056 367174
rect 156292 366938 156348 367174
rect 156000 366854 156348 366938
rect 156000 366618 156056 366854
rect 156292 366618 156348 366854
rect 156000 366586 156348 366618
rect 20952 363454 21300 363486
rect 20952 363218 21008 363454
rect 21244 363218 21300 363454
rect 20952 363134 21300 363218
rect 20952 362898 21008 363134
rect 21244 362898 21300 363134
rect 20952 362866 21300 362898
rect 155320 363454 155668 363486
rect 155320 363218 155376 363454
rect 155612 363218 155668 363454
rect 155320 363134 155668 363218
rect 155320 362898 155376 363134
rect 155612 362898 155668 363134
rect 155320 362866 155668 362898
rect 36056 349890 36116 350106
rect 37144 349890 37204 350106
rect 36056 349830 36186 349890
rect 37144 349830 37290 349890
rect 36126 347717 36186 349830
rect 36123 347716 36189 347717
rect 36123 347652 36124 347716
rect 36188 347652 36189 347716
rect 36123 347651 36189 347652
rect 37230 347309 37290 349830
rect 38232 349621 38292 350106
rect 39592 349890 39652 350106
rect 40544 349890 40604 350106
rect 39592 349830 39682 349890
rect 38229 349620 38295 349621
rect 38229 349556 38230 349620
rect 38294 349556 38295 349620
rect 38229 349555 38295 349556
rect 39622 347717 39682 349830
rect 40542 349830 40604 349890
rect 41768 349890 41828 350106
rect 43128 349890 43188 350106
rect 41768 349830 41890 349890
rect 39619 347716 39685 347717
rect 39619 347652 39620 347716
rect 39684 347652 39685 347716
rect 39619 347651 39685 347652
rect 37227 347308 37293 347309
rect 37227 347244 37228 347308
rect 37292 347244 37293 347308
rect 37227 347243 37293 347244
rect 40542 346493 40602 349830
rect 41830 346901 41890 349830
rect 43118 349830 43188 349890
rect 44216 349890 44276 350106
rect 45440 349890 45500 350106
rect 44216 349830 44282 349890
rect 43118 347717 43178 349830
rect 44222 347717 44282 349830
rect 45326 349830 45500 349890
rect 46528 349890 46588 350106
rect 47616 349890 47676 350106
rect 48296 349890 48356 350106
rect 48704 349890 48764 350106
rect 46528 349830 46674 349890
rect 45326 347717 45386 349830
rect 46614 347717 46674 349830
rect 47534 349830 47676 349890
rect 48270 349830 48356 349890
rect 48638 349830 48764 349890
rect 50064 349890 50124 350106
rect 50064 349830 50170 349890
rect 47534 347717 47594 349830
rect 43115 347716 43181 347717
rect 43115 347652 43116 347716
rect 43180 347652 43181 347716
rect 43115 347651 43181 347652
rect 44219 347716 44285 347717
rect 44219 347652 44220 347716
rect 44284 347652 44285 347716
rect 44219 347651 44285 347652
rect 45323 347716 45389 347717
rect 45323 347652 45324 347716
rect 45388 347652 45389 347716
rect 45323 347651 45389 347652
rect 46611 347716 46677 347717
rect 46611 347652 46612 347716
rect 46676 347652 46677 347716
rect 46611 347651 46677 347652
rect 47531 347716 47597 347717
rect 47531 347652 47532 347716
rect 47596 347652 47597 347716
rect 47531 347651 47597 347652
rect 48270 347581 48330 349830
rect 48638 347717 48698 349830
rect 50110 347717 50170 349830
rect 50744 349621 50804 350106
rect 51288 349890 51348 350106
rect 52376 349890 52436 350106
rect 53464 349890 53524 350106
rect 51214 349830 51348 349890
rect 52318 349830 52436 349890
rect 53422 349830 53524 349890
rect 53600 349890 53660 350106
rect 54552 349890 54612 350106
rect 55912 349890 55972 350106
rect 53600 349830 53666 349890
rect 50741 349620 50807 349621
rect 50741 349556 50742 349620
rect 50806 349556 50807 349620
rect 50741 349555 50807 349556
rect 51214 347717 51274 349830
rect 52318 347717 52378 349830
rect 53422 347717 53482 349830
rect 53606 349077 53666 349830
rect 54526 349830 54612 349890
rect 55814 349830 55972 349890
rect 53603 349076 53669 349077
rect 53603 349012 53604 349076
rect 53668 349012 53669 349076
rect 53603 349011 53669 349012
rect 48635 347716 48701 347717
rect 48635 347652 48636 347716
rect 48700 347652 48701 347716
rect 48635 347651 48701 347652
rect 50107 347716 50173 347717
rect 50107 347652 50108 347716
rect 50172 347652 50173 347716
rect 50107 347651 50173 347652
rect 51211 347716 51277 347717
rect 51211 347652 51212 347716
rect 51276 347652 51277 347716
rect 51211 347651 51277 347652
rect 52315 347716 52381 347717
rect 52315 347652 52316 347716
rect 52380 347652 52381 347716
rect 52315 347651 52381 347652
rect 53419 347716 53485 347717
rect 53419 347652 53420 347716
rect 53484 347652 53485 347716
rect 53419 347651 53485 347652
rect 48267 347580 48333 347581
rect 48267 347516 48268 347580
rect 48332 347516 48333 347580
rect 48267 347515 48333 347516
rect 41827 346900 41893 346901
rect 41827 346836 41828 346900
rect 41892 346836 41893 346900
rect 41827 346835 41893 346836
rect 54526 346765 54586 349830
rect 55814 347445 55874 349830
rect 56048 349621 56108 350106
rect 57000 349890 57060 350106
rect 58088 349890 58148 350106
rect 57000 349830 57162 349890
rect 58088 349830 58266 349890
rect 56045 349620 56111 349621
rect 56045 349556 56046 349620
rect 56110 349556 56111 349620
rect 56045 349555 56111 349556
rect 55811 347444 55877 347445
rect 55811 347380 55812 347444
rect 55876 347380 55877 347444
rect 55811 347379 55877 347380
rect 57102 347173 57162 349830
rect 58206 347445 58266 349830
rect 58496 349621 58556 350106
rect 59448 349890 59508 350106
rect 60672 349890 60732 350106
rect 59448 349830 59554 349890
rect 58493 349620 58559 349621
rect 58493 349556 58494 349620
rect 58558 349556 58559 349620
rect 58493 349555 58559 349556
rect 59494 347445 59554 349830
rect 60598 349830 60732 349890
rect 58203 347444 58269 347445
rect 58203 347380 58204 347444
rect 58268 347380 58269 347444
rect 58203 347379 58269 347380
rect 59491 347444 59557 347445
rect 59491 347380 59492 347444
rect 59556 347380 59557 347444
rect 59491 347379 59557 347380
rect 60598 347173 60658 349830
rect 61080 349621 61140 350106
rect 61760 349890 61820 350106
rect 61760 349830 61946 349890
rect 61077 349620 61143 349621
rect 61077 349556 61078 349620
rect 61142 349556 61143 349620
rect 61077 349555 61143 349556
rect 61886 349077 61946 349830
rect 62848 349621 62908 350106
rect 63528 349890 63588 350106
rect 63936 349890 63996 350106
rect 65296 349890 65356 350106
rect 65976 349890 66036 350106
rect 66384 349890 66444 350106
rect 67608 349890 67668 350106
rect 63528 349830 63602 349890
rect 62845 349620 62911 349621
rect 62845 349556 62846 349620
rect 62910 349556 62911 349620
rect 62845 349555 62911 349556
rect 61883 349076 61949 349077
rect 61883 349012 61884 349076
rect 61948 349012 61949 349076
rect 61883 349011 61949 349012
rect 63542 347717 63602 349830
rect 63910 349830 63996 349890
rect 65198 349830 65356 349890
rect 65934 349830 66036 349890
rect 66302 349830 66444 349890
rect 67590 349830 67668 349890
rect 68288 349890 68348 350106
rect 68288 349830 68386 349890
rect 63910 347717 63970 349830
rect 65198 347717 65258 349830
rect 65934 347717 65994 349830
rect 66302 347717 66362 349830
rect 67590 347717 67650 349830
rect 68326 349077 68386 349830
rect 68696 349621 68756 350106
rect 69784 349890 69844 350106
rect 71008 349890 71068 350106
rect 69784 349830 69858 349890
rect 68693 349620 68759 349621
rect 68693 349556 68694 349620
rect 68758 349556 68759 349620
rect 68693 349555 68759 349556
rect 68323 349076 68389 349077
rect 68323 349012 68324 349076
rect 68388 349012 68389 349076
rect 68323 349011 68389 349012
rect 63539 347716 63605 347717
rect 63539 347652 63540 347716
rect 63604 347652 63605 347716
rect 63539 347651 63605 347652
rect 63907 347716 63973 347717
rect 63907 347652 63908 347716
rect 63972 347652 63973 347716
rect 63907 347651 63973 347652
rect 65195 347716 65261 347717
rect 65195 347652 65196 347716
rect 65260 347652 65261 347716
rect 65195 347651 65261 347652
rect 65931 347716 65997 347717
rect 65931 347652 65932 347716
rect 65996 347652 65997 347716
rect 65931 347651 65997 347652
rect 66299 347716 66365 347717
rect 66299 347652 66300 347716
rect 66364 347652 66365 347716
rect 66299 347651 66365 347652
rect 67587 347716 67653 347717
rect 67587 347652 67588 347716
rect 67652 347652 67653 347716
rect 67587 347651 67653 347652
rect 69798 347173 69858 349830
rect 70902 349830 71068 349890
rect 71144 349890 71204 350106
rect 71144 349830 71330 349890
rect 70902 347445 70962 349830
rect 71270 347717 71330 349830
rect 72232 349621 72292 350106
rect 73320 349890 73380 350106
rect 73294 349830 73380 349890
rect 73592 349890 73652 350106
rect 74408 349890 74468 350106
rect 75768 349890 75828 350106
rect 73592 349830 73722 349890
rect 72229 349620 72295 349621
rect 72229 349556 72230 349620
rect 72294 349556 72295 349620
rect 72229 349555 72295 349556
rect 73294 347717 73354 349830
rect 73662 347717 73722 349830
rect 74398 349830 74468 349890
rect 75686 349830 75828 349890
rect 74398 348533 74458 349830
rect 74395 348532 74461 348533
rect 74395 348468 74396 348532
rect 74460 348468 74461 348532
rect 74395 348467 74461 348468
rect 75686 347717 75746 349830
rect 76040 349618 76100 350106
rect 76992 349618 77052 350106
rect 78080 349618 78140 350106
rect 78488 349618 78548 350106
rect 76040 349558 76114 349618
rect 76054 347717 76114 349558
rect 76974 349558 77052 349618
rect 78078 349558 78140 349618
rect 78446 349558 78548 349618
rect 79168 349618 79228 350106
rect 80936 349890 80996 350106
rect 83520 349890 83580 350106
rect 85968 349890 86028 350106
rect 88280 349890 88340 350106
rect 91000 349893 91060 350106
rect 93448 349893 93508 350106
rect 80936 349830 81082 349890
rect 83520 349830 83658 349890
rect 85968 349830 86050 349890
rect 79168 349558 79242 349618
rect 76974 347717 77034 349558
rect 78078 347717 78138 349558
rect 78446 349077 78506 349558
rect 78443 349076 78509 349077
rect 78443 349012 78444 349076
rect 78508 349012 78509 349076
rect 78443 349011 78509 349012
rect 79182 347717 79242 349558
rect 81022 347717 81082 349830
rect 83598 347717 83658 349830
rect 85990 349077 86050 349830
rect 88198 349830 88340 349890
rect 90997 349892 91063 349893
rect 88198 349077 88258 349830
rect 90997 349828 90998 349892
rect 91062 349828 91063 349892
rect 90997 349827 91063 349828
rect 93445 349892 93511 349893
rect 93445 349828 93446 349892
rect 93510 349828 93511 349892
rect 93445 349827 93511 349828
rect 95896 349618 95956 350106
rect 98480 349893 98540 350106
rect 98477 349892 98543 349893
rect 98477 349828 98478 349892
rect 98542 349828 98543 349892
rect 98477 349827 98543 349828
rect 100928 349618 100988 350106
rect 103512 349893 103572 350106
rect 103509 349892 103575 349893
rect 103509 349828 103510 349892
rect 103574 349828 103575 349892
rect 105960 349890 106020 350106
rect 108544 349890 108604 350106
rect 110992 349890 111052 350106
rect 113440 349890 113500 350106
rect 115888 349890 115948 350106
rect 105960 349830 106106 349890
rect 108544 349830 108682 349890
rect 110992 349830 111074 349890
rect 103509 349827 103575 349828
rect 95896 349558 95986 349618
rect 85987 349076 86053 349077
rect 85987 349012 85988 349076
rect 86052 349012 86053 349076
rect 85987 349011 86053 349012
rect 88195 349076 88261 349077
rect 88195 349012 88196 349076
rect 88260 349012 88261 349076
rect 88195 349011 88261 349012
rect 95926 347717 95986 349558
rect 100894 349558 100988 349618
rect 100894 347717 100954 349558
rect 106046 347717 106106 349830
rect 108622 347717 108682 349830
rect 111014 347717 111074 349830
rect 113406 349830 113500 349890
rect 115798 349830 115948 349890
rect 118472 349890 118532 350106
rect 120920 349890 120980 350106
rect 123368 349890 123428 350106
rect 125952 349890 126012 350106
rect 118472 349830 118618 349890
rect 120920 349830 121010 349890
rect 113406 347717 113466 349830
rect 115798 347717 115858 349830
rect 118558 347717 118618 349830
rect 120950 347717 121010 349830
rect 123342 349830 123428 349890
rect 125918 349830 126012 349890
rect 123342 347717 123402 349830
rect 125918 347717 125978 349830
rect 71267 347716 71333 347717
rect 71267 347652 71268 347716
rect 71332 347652 71333 347716
rect 71267 347651 71333 347652
rect 73291 347716 73357 347717
rect 73291 347652 73292 347716
rect 73356 347652 73357 347716
rect 73291 347651 73357 347652
rect 73659 347716 73725 347717
rect 73659 347652 73660 347716
rect 73724 347652 73725 347716
rect 73659 347651 73725 347652
rect 75683 347716 75749 347717
rect 75683 347652 75684 347716
rect 75748 347652 75749 347716
rect 75683 347651 75749 347652
rect 76051 347716 76117 347717
rect 76051 347652 76052 347716
rect 76116 347652 76117 347716
rect 76051 347651 76117 347652
rect 76971 347716 77037 347717
rect 76971 347652 76972 347716
rect 77036 347652 77037 347716
rect 76971 347651 77037 347652
rect 78075 347716 78141 347717
rect 78075 347652 78076 347716
rect 78140 347652 78141 347716
rect 78075 347651 78141 347652
rect 79179 347716 79245 347717
rect 79179 347652 79180 347716
rect 79244 347652 79245 347716
rect 79179 347651 79245 347652
rect 81019 347716 81085 347717
rect 81019 347652 81020 347716
rect 81084 347652 81085 347716
rect 81019 347651 81085 347652
rect 83595 347716 83661 347717
rect 83595 347652 83596 347716
rect 83660 347652 83661 347716
rect 83595 347651 83661 347652
rect 95923 347716 95989 347717
rect 95923 347652 95924 347716
rect 95988 347652 95989 347716
rect 95923 347651 95989 347652
rect 100891 347716 100957 347717
rect 100891 347652 100892 347716
rect 100956 347652 100957 347716
rect 100891 347651 100957 347652
rect 106043 347716 106109 347717
rect 106043 347652 106044 347716
rect 106108 347652 106109 347716
rect 106043 347651 106109 347652
rect 108619 347716 108685 347717
rect 108619 347652 108620 347716
rect 108684 347652 108685 347716
rect 108619 347651 108685 347652
rect 111011 347716 111077 347717
rect 111011 347652 111012 347716
rect 111076 347652 111077 347716
rect 111011 347651 111077 347652
rect 113403 347716 113469 347717
rect 113403 347652 113404 347716
rect 113468 347652 113469 347716
rect 113403 347651 113469 347652
rect 115795 347716 115861 347717
rect 115795 347652 115796 347716
rect 115860 347652 115861 347716
rect 115795 347651 115861 347652
rect 118555 347716 118621 347717
rect 118555 347652 118556 347716
rect 118620 347652 118621 347716
rect 118555 347651 118621 347652
rect 120947 347716 121013 347717
rect 120947 347652 120948 347716
rect 121012 347652 121013 347716
rect 120947 347651 121013 347652
rect 123339 347716 123405 347717
rect 123339 347652 123340 347716
rect 123404 347652 123405 347716
rect 123339 347651 123405 347652
rect 125915 347716 125981 347717
rect 125915 347652 125916 347716
rect 125980 347652 125981 347716
rect 125915 347651 125981 347652
rect 70899 347444 70965 347445
rect 70899 347380 70900 347444
rect 70964 347380 70965 347444
rect 70899 347379 70965 347380
rect 57099 347172 57165 347173
rect 57099 347108 57100 347172
rect 57164 347108 57165 347172
rect 57099 347107 57165 347108
rect 60595 347172 60661 347173
rect 60595 347108 60596 347172
rect 60660 347108 60661 347172
rect 60595 347107 60661 347108
rect 69795 347172 69861 347173
rect 69795 347108 69796 347172
rect 69860 347108 69861 347172
rect 69795 347107 69861 347108
rect 54523 346764 54589 346765
rect 54523 346700 54524 346764
rect 54588 346700 54589 346764
rect 54523 346699 54589 346700
rect 40539 346492 40605 346493
rect 40539 346428 40540 346492
rect 40604 346428 40605 346492
rect 40539 346427 40605 346428
rect 160674 342334 161294 377778
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 150939 335476 151005 335477
rect 150939 335412 150940 335476
rect 151004 335412 151005 335476
rect 150939 335411 151005 335412
rect 150942 333570 151002 335411
rect 150840 333510 151002 333570
rect 150840 333202 150900 333510
rect 20272 331174 20620 331206
rect 20272 330938 20328 331174
rect 20564 330938 20620 331174
rect 20272 330854 20620 330938
rect 20272 330618 20328 330854
rect 20564 330618 20620 330854
rect 20272 330586 20620 330618
rect 156000 331174 156348 331206
rect 156000 330938 156056 331174
rect 156292 330938 156348 331174
rect 156000 330854 156348 330938
rect 156000 330618 156056 330854
rect 156292 330618 156348 330854
rect 156000 330586 156348 330618
rect 20952 327454 21300 327486
rect 20952 327218 21008 327454
rect 21244 327218 21300 327454
rect 20952 327134 21300 327218
rect 20952 326898 21008 327134
rect 21244 326898 21300 327134
rect 20952 326866 21300 326898
rect 155320 327454 155668 327486
rect 155320 327218 155376 327454
rect 155612 327218 155668 327454
rect 155320 327134 155668 327218
rect 155320 326898 155376 327134
rect 155612 326898 155668 327134
rect 155320 326866 155668 326898
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 20272 295174 20620 295206
rect 20272 294938 20328 295174
rect 20564 294938 20620 295174
rect 20272 294854 20620 294938
rect 20272 294618 20328 294854
rect 20564 294618 20620 294854
rect 20272 294586 20620 294618
rect 156000 295174 156348 295206
rect 156000 294938 156056 295174
rect 156292 294938 156348 295174
rect 156000 294854 156348 294938
rect 156000 294618 156056 294854
rect 156292 294618 156348 294854
rect 156000 294586 156348 294618
rect 20952 291454 21300 291486
rect 20952 291218 21008 291454
rect 21244 291218 21300 291454
rect 20952 291134 21300 291218
rect 20952 290898 21008 291134
rect 21244 290898 21300 291134
rect 20952 290866 21300 290898
rect 155320 291454 155668 291486
rect 155320 291218 155376 291454
rect 155612 291218 155668 291454
rect 155320 291134 155668 291218
rect 155320 290898 155376 291134
rect 155612 290898 155668 291134
rect 155320 290866 155668 290898
rect 160674 270334 161294 305778
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 20272 259174 20620 259206
rect 20272 258938 20328 259174
rect 20564 258938 20620 259174
rect 20272 258854 20620 258938
rect 20272 258618 20328 258854
rect 20564 258618 20620 258854
rect 20272 258586 20620 258618
rect 156000 259174 156348 259206
rect 156000 258938 156056 259174
rect 156292 258938 156348 259174
rect 156000 258854 156348 258938
rect 156000 258618 156056 258854
rect 156292 258618 156348 258854
rect 156000 258586 156348 258618
rect 20952 255454 21300 255486
rect 20952 255218 21008 255454
rect 21244 255218 21300 255454
rect 20952 255134 21300 255218
rect 20952 254898 21008 255134
rect 21244 254898 21300 255134
rect 20952 254866 21300 254898
rect 155320 255454 155668 255486
rect 155320 255218 155376 255454
rect 155612 255218 155668 255454
rect 155320 255134 155668 255218
rect 155320 254898 155376 255134
rect 155612 254898 155668 255134
rect 155320 254866 155668 254898
rect 36056 249930 36116 250106
rect 37144 249930 37204 250106
rect 38232 249930 38292 250106
rect 35942 249870 36116 249930
rect 37046 249870 37204 249930
rect 38150 249870 38292 249930
rect 39592 249930 39652 250106
rect 40544 249930 40604 250106
rect 41768 249930 41828 250106
rect 43128 249930 43188 250106
rect 39592 249870 39682 249930
rect 35942 248301 36002 249870
rect 37046 248301 37106 249870
rect 35939 248300 36005 248301
rect 35939 248236 35940 248300
rect 36004 248236 36005 248300
rect 35939 248235 36005 248236
rect 37043 248300 37109 248301
rect 37043 248236 37044 248300
rect 37108 248236 37109 248300
rect 37043 248235 37109 248236
rect 38150 248165 38210 249870
rect 39622 248301 39682 249870
rect 40542 249870 40604 249930
rect 41646 249870 41828 249930
rect 43118 249870 43188 249930
rect 44216 249930 44276 250106
rect 45440 249930 45500 250106
rect 44216 249870 44282 249930
rect 39619 248300 39685 248301
rect 39619 248236 39620 248300
rect 39684 248236 39685 248300
rect 39619 248235 39685 248236
rect 40542 248165 40602 249870
rect 41646 248165 41706 249870
rect 43118 248165 43178 249870
rect 44222 248301 44282 249870
rect 45326 249870 45500 249930
rect 46528 249930 46588 250106
rect 47616 249930 47676 250106
rect 46528 249870 46674 249930
rect 44219 248300 44285 248301
rect 44219 248236 44220 248300
rect 44284 248236 44285 248300
rect 44219 248235 44285 248236
rect 45326 248165 45386 249870
rect 46614 248301 46674 249870
rect 47534 249870 47676 249930
rect 48296 249930 48356 250106
rect 48704 249930 48764 250106
rect 48296 249870 48514 249930
rect 46611 248300 46677 248301
rect 46611 248236 46612 248300
rect 46676 248236 46677 248300
rect 46611 248235 46677 248236
rect 47534 248165 47594 249870
rect 48454 248165 48514 249870
rect 48638 249870 48764 249930
rect 50064 249930 50124 250106
rect 50064 249870 50170 249930
rect 38147 248164 38213 248165
rect 38147 248100 38148 248164
rect 38212 248100 38213 248164
rect 38147 248099 38213 248100
rect 40539 248164 40605 248165
rect 40539 248100 40540 248164
rect 40604 248100 40605 248164
rect 40539 248099 40605 248100
rect 41643 248164 41709 248165
rect 41643 248100 41644 248164
rect 41708 248100 41709 248164
rect 41643 248099 41709 248100
rect 43115 248164 43181 248165
rect 43115 248100 43116 248164
rect 43180 248100 43181 248164
rect 43115 248099 43181 248100
rect 45323 248164 45389 248165
rect 45323 248100 45324 248164
rect 45388 248100 45389 248164
rect 45323 248099 45389 248100
rect 47531 248164 47597 248165
rect 47531 248100 47532 248164
rect 47596 248100 47597 248164
rect 47531 248099 47597 248100
rect 48451 248164 48517 248165
rect 48451 248100 48452 248164
rect 48516 248100 48517 248164
rect 48451 248099 48517 248100
rect 48638 247893 48698 249870
rect 50110 248301 50170 249870
rect 50744 249661 50804 250106
rect 51288 249930 51348 250106
rect 52376 249930 52436 250106
rect 53464 249930 53524 250106
rect 51288 249870 51458 249930
rect 50741 249660 50807 249661
rect 50741 249596 50742 249660
rect 50806 249596 50807 249660
rect 50741 249595 50807 249596
rect 50107 248300 50173 248301
rect 50107 248236 50108 248300
rect 50172 248236 50173 248300
rect 50107 248235 50173 248236
rect 48635 247892 48701 247893
rect 48635 247828 48636 247892
rect 48700 247828 48701 247892
rect 48635 247827 48701 247828
rect 51398 247485 51458 249870
rect 52318 249870 52436 249930
rect 53422 249870 53524 249930
rect 51395 247484 51461 247485
rect 51395 247420 51396 247484
rect 51460 247420 51461 247484
rect 51395 247419 51461 247420
rect 52318 247077 52378 249870
rect 53422 247349 53482 249870
rect 53600 249661 53660 250106
rect 54552 249930 54612 250106
rect 55912 249930 55972 250106
rect 54526 249870 54612 249930
rect 55814 249870 55972 249930
rect 53597 249660 53663 249661
rect 53597 249596 53598 249660
rect 53662 249596 53663 249660
rect 53597 249595 53663 249596
rect 53419 247348 53485 247349
rect 53419 247284 53420 247348
rect 53484 247284 53485 247348
rect 53419 247283 53485 247284
rect 54526 247077 54586 249870
rect 55814 247077 55874 249870
rect 56048 249661 56108 250106
rect 57000 249930 57060 250106
rect 58088 249930 58148 250106
rect 57000 249870 57162 249930
rect 56045 249660 56111 249661
rect 56045 249596 56046 249660
rect 56110 249596 56111 249660
rect 56045 249595 56111 249596
rect 57102 247077 57162 249870
rect 58022 249870 58148 249930
rect 58022 247893 58082 249870
rect 58496 249661 58556 250106
rect 59448 249930 59508 250106
rect 60672 249930 60732 250106
rect 59448 249870 59554 249930
rect 58493 249660 58559 249661
rect 58493 249596 58494 249660
rect 58558 249596 58559 249660
rect 58493 249595 58559 249596
rect 59494 247893 59554 249870
rect 60598 249870 60732 249930
rect 61080 249930 61140 250106
rect 61760 249930 61820 250106
rect 62848 249930 62908 250106
rect 61080 249870 61210 249930
rect 60598 248029 60658 249870
rect 61150 248301 61210 249870
rect 61702 249870 61820 249930
rect 62806 249870 62908 249930
rect 63528 249930 63588 250106
rect 63936 249930 63996 250106
rect 65296 249930 65356 250106
rect 65976 249930 66036 250106
rect 66384 249930 66444 250106
rect 63528 249870 63602 249930
rect 61702 248301 61762 249870
rect 62806 248301 62866 249870
rect 63542 248301 63602 249870
rect 63910 249870 63996 249930
rect 65198 249870 65356 249930
rect 65934 249870 66036 249930
rect 66302 249870 66444 249930
rect 67608 249930 67668 250106
rect 68288 249930 68348 250106
rect 68696 249930 68756 250106
rect 67608 249870 67834 249930
rect 68288 249870 68386 249930
rect 61147 248300 61213 248301
rect 61147 248236 61148 248300
rect 61212 248236 61213 248300
rect 61147 248235 61213 248236
rect 61699 248300 61765 248301
rect 61699 248236 61700 248300
rect 61764 248236 61765 248300
rect 61699 248235 61765 248236
rect 62803 248300 62869 248301
rect 62803 248236 62804 248300
rect 62868 248236 62869 248300
rect 62803 248235 62869 248236
rect 63539 248300 63605 248301
rect 63539 248236 63540 248300
rect 63604 248236 63605 248300
rect 63539 248235 63605 248236
rect 63910 248029 63970 249870
rect 65198 248301 65258 249870
rect 65934 248301 65994 249870
rect 65195 248300 65261 248301
rect 65195 248236 65196 248300
rect 65260 248236 65261 248300
rect 65195 248235 65261 248236
rect 65931 248300 65997 248301
rect 65931 248236 65932 248300
rect 65996 248236 65997 248300
rect 65931 248235 65997 248236
rect 60595 248028 60661 248029
rect 60595 247964 60596 248028
rect 60660 247964 60661 248028
rect 60595 247963 60661 247964
rect 63907 248028 63973 248029
rect 63907 247964 63908 248028
rect 63972 247964 63973 248028
rect 63907 247963 63973 247964
rect 66302 247893 66362 249870
rect 67774 247893 67834 249870
rect 68326 247893 68386 249870
rect 68694 249870 68756 249930
rect 69784 249930 69844 250106
rect 71008 249930 71068 250106
rect 69784 249870 69858 249930
rect 68694 248301 68754 249870
rect 68691 248300 68757 248301
rect 68691 248236 68692 248300
rect 68756 248236 68757 248300
rect 68691 248235 68757 248236
rect 58019 247892 58085 247893
rect 58019 247828 58020 247892
rect 58084 247828 58085 247892
rect 58019 247827 58085 247828
rect 59491 247892 59557 247893
rect 59491 247828 59492 247892
rect 59556 247828 59557 247892
rect 59491 247827 59557 247828
rect 66299 247892 66365 247893
rect 66299 247828 66300 247892
rect 66364 247828 66365 247892
rect 66299 247827 66365 247828
rect 67771 247892 67837 247893
rect 67771 247828 67772 247892
rect 67836 247828 67837 247892
rect 67771 247827 67837 247828
rect 68323 247892 68389 247893
rect 68323 247828 68324 247892
rect 68388 247828 68389 247892
rect 68323 247827 68389 247828
rect 69798 247485 69858 249870
rect 70902 249870 71068 249930
rect 71144 249930 71204 250106
rect 72232 249930 72292 250106
rect 73320 249930 73380 250106
rect 71144 249870 71330 249930
rect 70902 248301 70962 249870
rect 70899 248300 70965 248301
rect 70899 248236 70900 248300
rect 70964 248236 70965 248300
rect 70899 248235 70965 248236
rect 69795 247484 69861 247485
rect 69795 247420 69796 247484
rect 69860 247420 69861 247484
rect 69795 247419 69861 247420
rect 71270 247349 71330 249870
rect 72190 249870 72292 249930
rect 73294 249870 73380 249930
rect 73592 249930 73652 250106
rect 74408 249930 74468 250106
rect 75768 249930 75828 250106
rect 73592 249870 73722 249930
rect 72190 247621 72250 249870
rect 72187 247620 72253 247621
rect 72187 247556 72188 247620
rect 72252 247556 72253 247620
rect 72187 247555 72253 247556
rect 71267 247348 71333 247349
rect 71267 247284 71268 247348
rect 71332 247284 71333 247348
rect 71267 247283 71333 247284
rect 73294 247213 73354 249870
rect 73662 248301 73722 249870
rect 74398 249870 74468 249930
rect 75686 249870 75828 249930
rect 76040 249930 76100 250106
rect 76992 249930 77052 250106
rect 78080 249930 78140 250106
rect 78488 249930 78548 250106
rect 76040 249870 76114 249930
rect 73659 248300 73725 248301
rect 73659 248236 73660 248300
rect 73724 248236 73725 248300
rect 73659 248235 73725 248236
rect 74398 247349 74458 249870
rect 75686 247757 75746 249870
rect 76054 247893 76114 249870
rect 76974 249870 77052 249930
rect 78078 249870 78140 249930
rect 78446 249870 78548 249930
rect 79168 249930 79228 250106
rect 80936 249930 80996 250106
rect 83520 249930 83580 250106
rect 85968 249930 86028 250106
rect 88280 249930 88340 250106
rect 91000 249930 91060 250106
rect 79168 249870 79242 249930
rect 80936 249870 81082 249930
rect 83520 249870 83658 249930
rect 85968 249870 86050 249930
rect 76051 247892 76117 247893
rect 76051 247828 76052 247892
rect 76116 247828 76117 247892
rect 76051 247827 76117 247828
rect 76974 247757 77034 249870
rect 78078 248301 78138 249870
rect 78446 248301 78506 249870
rect 78075 248300 78141 248301
rect 78075 248236 78076 248300
rect 78140 248236 78141 248300
rect 78075 248235 78141 248236
rect 78443 248300 78509 248301
rect 78443 248236 78444 248300
rect 78508 248236 78509 248300
rect 78443 248235 78509 248236
rect 79182 248029 79242 249870
rect 81022 248029 81082 249870
rect 83598 248301 83658 249870
rect 83595 248300 83661 248301
rect 83595 248236 83596 248300
rect 83660 248236 83661 248300
rect 83595 248235 83661 248236
rect 85990 248029 86050 249870
rect 88198 249870 88340 249930
rect 90958 249870 91060 249930
rect 88198 248029 88258 249870
rect 90958 248029 91018 249870
rect 93448 249797 93508 250106
rect 95896 249797 95956 250106
rect 98480 249797 98540 250106
rect 93445 249796 93511 249797
rect 93445 249732 93446 249796
rect 93510 249732 93511 249796
rect 93445 249731 93511 249732
rect 95893 249796 95959 249797
rect 95893 249732 95894 249796
rect 95958 249732 95959 249796
rect 95893 249731 95959 249732
rect 98477 249796 98543 249797
rect 98477 249732 98478 249796
rect 98542 249732 98543 249796
rect 100928 249794 100988 250106
rect 103512 249797 103572 250106
rect 105960 249797 106020 250106
rect 108544 249797 108604 250106
rect 110992 249797 111052 250106
rect 98477 249731 98543 249732
rect 100894 249734 100988 249794
rect 103509 249796 103575 249797
rect 100894 248029 100954 249734
rect 103509 249732 103510 249796
rect 103574 249732 103575 249796
rect 103509 249731 103575 249732
rect 105957 249796 106023 249797
rect 105957 249732 105958 249796
rect 106022 249732 106023 249796
rect 105957 249731 106023 249732
rect 108541 249796 108607 249797
rect 108541 249732 108542 249796
rect 108606 249732 108607 249796
rect 108541 249731 108607 249732
rect 110989 249796 111055 249797
rect 110989 249732 110990 249796
rect 111054 249732 111055 249796
rect 110989 249731 111055 249732
rect 113440 249661 113500 250106
rect 115888 249661 115948 250106
rect 118472 249930 118532 250106
rect 118472 249870 118618 249930
rect 113437 249660 113503 249661
rect 113437 249596 113438 249660
rect 113502 249596 113503 249660
rect 113437 249595 113503 249596
rect 115885 249660 115951 249661
rect 115885 249596 115886 249660
rect 115950 249596 115951 249660
rect 115885 249595 115951 249596
rect 118558 248029 118618 249870
rect 120920 249661 120980 250106
rect 123368 249930 123428 250106
rect 125952 249930 126012 250106
rect 123342 249870 123428 249930
rect 125918 249870 126012 249930
rect 120917 249660 120983 249661
rect 120917 249596 120918 249660
rect 120982 249596 120983 249660
rect 120917 249595 120983 249596
rect 79179 248028 79245 248029
rect 79179 247964 79180 248028
rect 79244 247964 79245 248028
rect 79179 247963 79245 247964
rect 81019 248028 81085 248029
rect 81019 247964 81020 248028
rect 81084 247964 81085 248028
rect 81019 247963 81085 247964
rect 85987 248028 86053 248029
rect 85987 247964 85988 248028
rect 86052 247964 86053 248028
rect 85987 247963 86053 247964
rect 88195 248028 88261 248029
rect 88195 247964 88196 248028
rect 88260 247964 88261 248028
rect 88195 247963 88261 247964
rect 90955 248028 91021 248029
rect 90955 247964 90956 248028
rect 91020 247964 91021 248028
rect 90955 247963 91021 247964
rect 100891 248028 100957 248029
rect 100891 247964 100892 248028
rect 100956 247964 100957 248028
rect 100891 247963 100957 247964
rect 118555 248028 118621 248029
rect 118555 247964 118556 248028
rect 118620 247964 118621 248028
rect 118555 247963 118621 247964
rect 123342 247893 123402 249870
rect 125918 248301 125978 249870
rect 125915 248300 125981 248301
rect 125915 248236 125916 248300
rect 125980 248236 125981 248300
rect 125915 248235 125981 248236
rect 123339 247892 123405 247893
rect 123339 247828 123340 247892
rect 123404 247828 123405 247892
rect 123339 247827 123405 247828
rect 75683 247756 75749 247757
rect 75683 247692 75684 247756
rect 75748 247692 75749 247756
rect 75683 247691 75749 247692
rect 76971 247756 77037 247757
rect 76971 247692 76972 247756
rect 77036 247692 77037 247756
rect 76971 247691 77037 247692
rect 74395 247348 74461 247349
rect 74395 247284 74396 247348
rect 74460 247284 74461 247348
rect 74395 247283 74461 247284
rect 73291 247212 73357 247213
rect 73291 247148 73292 247212
rect 73356 247148 73357 247212
rect 73291 247147 73357 247148
rect 52315 247076 52381 247077
rect 52315 247012 52316 247076
rect 52380 247012 52381 247076
rect 52315 247011 52381 247012
rect 54523 247076 54589 247077
rect 54523 247012 54524 247076
rect 54588 247012 54589 247076
rect 54523 247011 54589 247012
rect 55811 247076 55877 247077
rect 55811 247012 55812 247076
rect 55876 247012 55877 247076
rect 55811 247011 55877 247012
rect 57099 247076 57165 247077
rect 57099 247012 57100 247076
rect 57164 247012 57165 247076
rect 57099 247011 57165 247012
rect 150755 234700 150821 234701
rect 150755 234636 150756 234700
rect 150820 234636 150821 234700
rect 150755 234635 150821 234636
rect 150758 233610 150818 234635
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 150758 233550 150900 233610
rect 150840 233240 150900 233550
rect 20272 223174 20620 223206
rect 20272 222938 20328 223174
rect 20564 222938 20620 223174
rect 20272 222854 20620 222938
rect 20272 222618 20328 222854
rect 20564 222618 20620 222854
rect 20272 222586 20620 222618
rect 156000 223174 156348 223206
rect 156000 222938 156056 223174
rect 156292 222938 156348 223174
rect 156000 222854 156348 222938
rect 156000 222618 156056 222854
rect 156292 222618 156348 222854
rect 156000 222586 156348 222618
rect 20952 219454 21300 219486
rect 20952 219218 21008 219454
rect 21244 219218 21300 219454
rect 20952 219134 21300 219218
rect 20952 218898 21008 219134
rect 21244 218898 21300 219134
rect 20952 218866 21300 218898
rect 155320 219454 155668 219486
rect 155320 219218 155376 219454
rect 155612 219218 155668 219454
rect 155320 219134 155668 219218
rect 155320 218898 155376 219134
rect 155612 218898 155668 219134
rect 155320 218866 155668 218898
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 20272 187174 20620 187206
rect 20272 186938 20328 187174
rect 20564 186938 20620 187174
rect 20272 186854 20620 186938
rect 20272 186618 20328 186854
rect 20564 186618 20620 186854
rect 20272 186586 20620 186618
rect 156000 187174 156348 187206
rect 156000 186938 156056 187174
rect 156292 186938 156348 187174
rect 156000 186854 156348 186938
rect 156000 186618 156056 186854
rect 156292 186618 156348 186854
rect 156000 186586 156348 186618
rect 20952 183454 21300 183486
rect 20952 183218 21008 183454
rect 21244 183218 21300 183454
rect 20952 183134 21300 183218
rect 20952 182898 21008 183134
rect 21244 182898 21300 183134
rect 20952 182866 21300 182898
rect 155320 183454 155668 183486
rect 155320 183218 155376 183454
rect 155612 183218 155668 183454
rect 155320 183134 155668 183218
rect 155320 182898 155376 183134
rect 155612 182898 155668 183134
rect 155320 182866 155668 182898
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 20272 151174 20620 151206
rect 20272 150938 20328 151174
rect 20564 150938 20620 151174
rect 20272 150854 20620 150938
rect 20272 150618 20328 150854
rect 20564 150618 20620 150854
rect 20272 150586 20620 150618
rect 156000 151174 156348 151206
rect 156000 150938 156056 151174
rect 156292 150938 156348 151174
rect 156000 150854 156348 150938
rect 156000 150618 156056 150854
rect 156292 150618 156348 150854
rect 156000 150586 156348 150618
rect 36056 149290 36116 150106
rect 37144 149290 37204 150106
rect 38232 149290 38292 150106
rect 35942 149230 36116 149290
rect 37046 149230 37204 149290
rect 38150 149230 38292 149290
rect 39592 149290 39652 150106
rect 40544 149290 40604 150106
rect 39592 149230 39682 149290
rect 35942 147661 36002 149230
rect 37046 147661 37106 149230
rect 38150 147661 38210 149230
rect 39622 147661 39682 149230
rect 40542 149230 40604 149290
rect 41768 149290 41828 150106
rect 43128 149290 43188 150106
rect 41768 149230 41890 149290
rect 35939 147660 36005 147661
rect 35939 147596 35940 147660
rect 36004 147596 36005 147660
rect 35939 147595 36005 147596
rect 37043 147660 37109 147661
rect 37043 147596 37044 147660
rect 37108 147596 37109 147660
rect 37043 147595 37109 147596
rect 38147 147660 38213 147661
rect 38147 147596 38148 147660
rect 38212 147596 38213 147660
rect 38147 147595 38213 147596
rect 39619 147660 39685 147661
rect 39619 147596 39620 147660
rect 39684 147596 39685 147660
rect 39619 147595 39685 147596
rect 40542 147389 40602 149230
rect 41830 147525 41890 149230
rect 43118 149230 43188 149290
rect 44216 149290 44276 150106
rect 45440 149290 45500 150106
rect 44216 149230 44282 149290
rect 43118 147661 43178 149230
rect 44222 147661 44282 149230
rect 45326 149230 45500 149290
rect 46528 149290 46588 150106
rect 47616 149290 47676 150106
rect 48296 149565 48356 150106
rect 48293 149564 48359 149565
rect 48293 149500 48294 149564
rect 48358 149500 48359 149564
rect 48293 149499 48359 149500
rect 48704 149290 48764 150106
rect 46528 149230 46674 149290
rect 47616 149230 47778 149290
rect 45326 147661 45386 149230
rect 46614 147661 46674 149230
rect 47718 147661 47778 149230
rect 48638 149230 48764 149290
rect 50064 149290 50124 150106
rect 50744 149565 50804 150106
rect 50741 149564 50807 149565
rect 50741 149500 50742 149564
rect 50806 149500 50807 149564
rect 50741 149499 50807 149500
rect 51288 149290 51348 150106
rect 52376 149290 52436 150106
rect 53464 149290 53524 150106
rect 50064 149230 50170 149290
rect 51288 149230 51458 149290
rect 48638 147661 48698 149230
rect 50110 147661 50170 149230
rect 51398 147661 51458 149230
rect 52318 149230 52436 149290
rect 53422 149230 53524 149290
rect 53600 149290 53660 150106
rect 54552 149290 54612 150106
rect 53600 149230 53666 149290
rect 52318 147661 52378 149230
rect 53422 147661 53482 149230
rect 53606 149021 53666 149230
rect 54526 149230 54612 149290
rect 55912 149290 55972 150106
rect 56048 149565 56108 150106
rect 56045 149564 56111 149565
rect 56045 149500 56046 149564
rect 56110 149500 56111 149564
rect 56045 149499 56111 149500
rect 57000 149290 57060 150106
rect 58088 149290 58148 150106
rect 58496 149565 58556 150106
rect 58493 149564 58559 149565
rect 58493 149500 58494 149564
rect 58558 149500 58559 149564
rect 58493 149499 58559 149500
rect 55912 149230 56058 149290
rect 53603 149020 53669 149021
rect 53603 148956 53604 149020
rect 53668 148956 53669 149020
rect 53603 148955 53669 148956
rect 54526 147661 54586 149230
rect 55998 147661 56058 149230
rect 56918 149230 57060 149290
rect 58022 149230 58148 149290
rect 59448 149290 59508 150106
rect 60672 149565 60732 150106
rect 60669 149564 60735 149565
rect 60669 149500 60670 149564
rect 60734 149500 60735 149564
rect 61080 149562 61140 150106
rect 61760 149562 61820 150106
rect 62848 149562 62908 150106
rect 61080 149502 61210 149562
rect 60669 149499 60735 149500
rect 59448 149230 59554 149290
rect 43115 147660 43181 147661
rect 43115 147596 43116 147660
rect 43180 147596 43181 147660
rect 43115 147595 43181 147596
rect 44219 147660 44285 147661
rect 44219 147596 44220 147660
rect 44284 147596 44285 147660
rect 44219 147595 44285 147596
rect 45323 147660 45389 147661
rect 45323 147596 45324 147660
rect 45388 147596 45389 147660
rect 45323 147595 45389 147596
rect 46611 147660 46677 147661
rect 46611 147596 46612 147660
rect 46676 147596 46677 147660
rect 46611 147595 46677 147596
rect 47715 147660 47781 147661
rect 47715 147596 47716 147660
rect 47780 147596 47781 147660
rect 47715 147595 47781 147596
rect 48635 147660 48701 147661
rect 48635 147596 48636 147660
rect 48700 147596 48701 147660
rect 48635 147595 48701 147596
rect 50107 147660 50173 147661
rect 50107 147596 50108 147660
rect 50172 147596 50173 147660
rect 50107 147595 50173 147596
rect 51395 147660 51461 147661
rect 51395 147596 51396 147660
rect 51460 147596 51461 147660
rect 51395 147595 51461 147596
rect 52315 147660 52381 147661
rect 52315 147596 52316 147660
rect 52380 147596 52381 147660
rect 52315 147595 52381 147596
rect 53419 147660 53485 147661
rect 53419 147596 53420 147660
rect 53484 147596 53485 147660
rect 53419 147595 53485 147596
rect 54523 147660 54589 147661
rect 54523 147596 54524 147660
rect 54588 147596 54589 147660
rect 54523 147595 54589 147596
rect 55995 147660 56061 147661
rect 55995 147596 55996 147660
rect 56060 147596 56061 147660
rect 55995 147595 56061 147596
rect 41827 147524 41893 147525
rect 41827 147460 41828 147524
rect 41892 147460 41893 147524
rect 41827 147459 41893 147460
rect 40539 147388 40605 147389
rect 40539 147324 40540 147388
rect 40604 147324 40605 147388
rect 40539 147323 40605 147324
rect 56918 147253 56978 149230
rect 58022 147661 58082 149230
rect 59494 147661 59554 149230
rect 58019 147660 58085 147661
rect 58019 147596 58020 147660
rect 58084 147596 58085 147660
rect 58019 147595 58085 147596
rect 59491 147660 59557 147661
rect 59491 147596 59492 147660
rect 59556 147596 59557 147660
rect 59491 147595 59557 147596
rect 61150 147389 61210 149502
rect 61702 149502 61820 149562
rect 62806 149502 62908 149562
rect 63528 149562 63588 150106
rect 63936 149562 63996 150106
rect 65296 149562 65356 150106
rect 63528 149502 63602 149562
rect 61702 147661 61762 149502
rect 62806 147661 62866 149502
rect 63542 147661 63602 149502
rect 63910 149502 63996 149562
rect 65198 149502 65356 149562
rect 65976 149562 66036 150106
rect 66384 149562 66444 150106
rect 67608 149562 67668 150106
rect 68288 149562 68348 150106
rect 68696 149562 68756 150106
rect 65976 149502 66178 149562
rect 63910 147661 63970 149502
rect 65198 147661 65258 149502
rect 66118 147661 66178 149502
rect 66302 149502 66444 149562
rect 67590 149502 67668 149562
rect 68142 149502 68348 149562
rect 68694 149502 68756 149562
rect 69784 149562 69844 150106
rect 71008 149565 71068 150106
rect 71005 149564 71071 149565
rect 69784 149502 69858 149562
rect 66302 147661 66362 149502
rect 67590 147661 67650 149502
rect 68142 147661 68202 149502
rect 68694 147661 68754 149502
rect 69798 147661 69858 149502
rect 71005 149500 71006 149564
rect 71070 149500 71071 149564
rect 71005 149499 71071 149500
rect 71144 149290 71204 150106
rect 72232 149290 72292 150106
rect 73320 149290 73380 150106
rect 73592 149565 73652 150106
rect 73589 149564 73655 149565
rect 73589 149500 73590 149564
rect 73654 149500 73655 149564
rect 73589 149499 73655 149500
rect 74408 149290 74468 150106
rect 75768 149290 75828 150106
rect 71086 149230 71204 149290
rect 72190 149230 72292 149290
rect 73294 149230 73380 149290
rect 74398 149230 74468 149290
rect 75686 149230 75828 149290
rect 76040 149290 76100 150106
rect 76992 149290 77052 150106
rect 78080 149290 78140 150106
rect 78488 149290 78548 150106
rect 76040 149230 76114 149290
rect 61699 147660 61765 147661
rect 61699 147596 61700 147660
rect 61764 147596 61765 147660
rect 61699 147595 61765 147596
rect 62803 147660 62869 147661
rect 62803 147596 62804 147660
rect 62868 147596 62869 147660
rect 62803 147595 62869 147596
rect 63539 147660 63605 147661
rect 63539 147596 63540 147660
rect 63604 147596 63605 147660
rect 63539 147595 63605 147596
rect 63907 147660 63973 147661
rect 63907 147596 63908 147660
rect 63972 147596 63973 147660
rect 63907 147595 63973 147596
rect 65195 147660 65261 147661
rect 65195 147596 65196 147660
rect 65260 147596 65261 147660
rect 65195 147595 65261 147596
rect 66115 147660 66181 147661
rect 66115 147596 66116 147660
rect 66180 147596 66181 147660
rect 66115 147595 66181 147596
rect 66299 147660 66365 147661
rect 66299 147596 66300 147660
rect 66364 147596 66365 147660
rect 66299 147595 66365 147596
rect 67587 147660 67653 147661
rect 67587 147596 67588 147660
rect 67652 147596 67653 147660
rect 67587 147595 67653 147596
rect 68139 147660 68205 147661
rect 68139 147596 68140 147660
rect 68204 147596 68205 147660
rect 68139 147595 68205 147596
rect 68691 147660 68757 147661
rect 68691 147596 68692 147660
rect 68756 147596 68757 147660
rect 68691 147595 68757 147596
rect 69795 147660 69861 147661
rect 69795 147596 69796 147660
rect 69860 147596 69861 147660
rect 69795 147595 69861 147596
rect 61147 147388 61213 147389
rect 61147 147324 61148 147388
rect 61212 147324 61213 147388
rect 61147 147323 61213 147324
rect 71086 147253 71146 149230
rect 72190 147661 72250 149230
rect 73294 147661 73354 149230
rect 74398 147661 74458 149230
rect 75686 147661 75746 149230
rect 76054 149021 76114 149230
rect 76974 149230 77052 149290
rect 78078 149230 78140 149290
rect 78446 149230 78548 149290
rect 79168 149290 79228 150106
rect 80936 149290 80996 150106
rect 83520 149565 83580 150106
rect 83517 149564 83583 149565
rect 83517 149500 83518 149564
rect 83582 149500 83583 149564
rect 83517 149499 83583 149500
rect 85968 149290 86028 150106
rect 88280 149290 88340 150106
rect 91000 149290 91060 150106
rect 93448 149565 93508 150106
rect 93445 149564 93511 149565
rect 93445 149500 93446 149564
rect 93510 149500 93511 149564
rect 93445 149499 93511 149500
rect 79168 149230 79242 149290
rect 80936 149230 81082 149290
rect 85968 149230 86050 149290
rect 76051 149020 76117 149021
rect 76051 148956 76052 149020
rect 76116 148956 76117 149020
rect 76051 148955 76117 148956
rect 76974 147661 77034 149230
rect 78078 147661 78138 149230
rect 78446 147661 78506 149230
rect 79182 147661 79242 149230
rect 81022 147661 81082 149230
rect 85990 149021 86050 149230
rect 88198 149230 88340 149290
rect 90958 149230 91060 149290
rect 95896 149290 95956 150106
rect 98480 149565 98540 150106
rect 98477 149564 98543 149565
rect 98477 149500 98478 149564
rect 98542 149500 98543 149564
rect 98477 149499 98543 149500
rect 100928 149290 100988 150106
rect 103512 149565 103572 150106
rect 103509 149564 103575 149565
rect 103509 149500 103510 149564
rect 103574 149500 103575 149564
rect 103509 149499 103575 149500
rect 95896 149230 95986 149290
rect 85987 149020 86053 149021
rect 85987 148956 85988 149020
rect 86052 148956 86053 149020
rect 85987 148955 86053 148956
rect 88198 147661 88258 149230
rect 90958 147661 91018 149230
rect 95926 147661 95986 149230
rect 100894 149230 100988 149290
rect 105960 149290 106020 150106
rect 108544 149290 108604 150106
rect 110992 149562 111052 150106
rect 113440 149565 113500 150106
rect 115888 149565 115948 150106
rect 113437 149564 113503 149565
rect 110992 149502 111074 149562
rect 105960 149230 106106 149290
rect 108544 149230 108682 149290
rect 100894 147661 100954 149230
rect 106046 147661 106106 149230
rect 108622 147661 108682 149230
rect 111014 147661 111074 149502
rect 113437 149500 113438 149564
rect 113502 149500 113503 149564
rect 113437 149499 113503 149500
rect 115885 149564 115951 149565
rect 115885 149500 115886 149564
rect 115950 149500 115951 149564
rect 115885 149499 115951 149500
rect 118472 149290 118532 150106
rect 120920 149565 120980 150106
rect 120917 149564 120983 149565
rect 120917 149500 120918 149564
rect 120982 149500 120983 149564
rect 120917 149499 120983 149500
rect 123368 149290 123428 150106
rect 125952 149290 126012 150106
rect 118472 149230 118618 149290
rect 72187 147660 72253 147661
rect 72187 147596 72188 147660
rect 72252 147596 72253 147660
rect 72187 147595 72253 147596
rect 73291 147660 73357 147661
rect 73291 147596 73292 147660
rect 73356 147596 73357 147660
rect 73291 147595 73357 147596
rect 74395 147660 74461 147661
rect 74395 147596 74396 147660
rect 74460 147596 74461 147660
rect 74395 147595 74461 147596
rect 75683 147660 75749 147661
rect 75683 147596 75684 147660
rect 75748 147596 75749 147660
rect 75683 147595 75749 147596
rect 76971 147660 77037 147661
rect 76971 147596 76972 147660
rect 77036 147596 77037 147660
rect 76971 147595 77037 147596
rect 78075 147660 78141 147661
rect 78075 147596 78076 147660
rect 78140 147596 78141 147660
rect 78075 147595 78141 147596
rect 78443 147660 78509 147661
rect 78443 147596 78444 147660
rect 78508 147596 78509 147660
rect 78443 147595 78509 147596
rect 79179 147660 79245 147661
rect 79179 147596 79180 147660
rect 79244 147596 79245 147660
rect 79179 147595 79245 147596
rect 81019 147660 81085 147661
rect 81019 147596 81020 147660
rect 81084 147596 81085 147660
rect 81019 147595 81085 147596
rect 88195 147660 88261 147661
rect 88195 147596 88196 147660
rect 88260 147596 88261 147660
rect 88195 147595 88261 147596
rect 90955 147660 91021 147661
rect 90955 147596 90956 147660
rect 91020 147596 91021 147660
rect 90955 147595 91021 147596
rect 95923 147660 95989 147661
rect 95923 147596 95924 147660
rect 95988 147596 95989 147660
rect 95923 147595 95989 147596
rect 100891 147660 100957 147661
rect 100891 147596 100892 147660
rect 100956 147596 100957 147660
rect 100891 147595 100957 147596
rect 106043 147660 106109 147661
rect 106043 147596 106044 147660
rect 106108 147596 106109 147660
rect 106043 147595 106109 147596
rect 108619 147660 108685 147661
rect 108619 147596 108620 147660
rect 108684 147596 108685 147660
rect 108619 147595 108685 147596
rect 111011 147660 111077 147661
rect 111011 147596 111012 147660
rect 111076 147596 111077 147660
rect 111011 147595 111077 147596
rect 118558 147525 118618 149230
rect 123342 149230 123428 149290
rect 125918 149230 126012 149290
rect 123342 149021 123402 149230
rect 123339 149020 123405 149021
rect 123339 148956 123340 149020
rect 123404 148956 123405 149020
rect 123339 148955 123405 148956
rect 125918 148885 125978 149230
rect 125915 148884 125981 148885
rect 125915 148820 125916 148884
rect 125980 148820 125981 148884
rect 125915 148819 125981 148820
rect 118555 147524 118621 147525
rect 118555 147460 118556 147524
rect 118620 147460 118621 147524
rect 118555 147459 118621 147460
rect 56915 147252 56981 147253
rect 56915 147188 56916 147252
rect 56980 147188 56981 147252
rect 56915 147187 56981 147188
rect 71083 147252 71149 147253
rect 71083 147188 71084 147252
rect 71148 147188 71149 147252
rect 71083 147187 71149 147188
rect 151123 135828 151189 135829
rect 151123 135764 151124 135828
rect 151188 135764 151189 135828
rect 151123 135763 151189 135764
rect 151126 133310 151186 135763
rect 150870 133250 151186 133310
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 20272 115174 20620 115206
rect 20272 114938 20328 115174
rect 20564 114938 20620 115174
rect 20272 114854 20620 114938
rect 20272 114618 20328 114854
rect 20564 114618 20620 114854
rect 20272 114586 20620 114618
rect 156000 115174 156348 115206
rect 156000 114938 156056 115174
rect 156292 114938 156348 115174
rect 156000 114854 156348 114938
rect 156000 114618 156056 114854
rect 156292 114618 156348 114854
rect 156000 114586 156348 114618
rect 20952 111454 21300 111486
rect 20952 111218 21008 111454
rect 21244 111218 21300 111454
rect 20952 111134 21300 111218
rect 20952 110898 21008 111134
rect 21244 110898 21300 111134
rect 20952 110866 21300 110898
rect 155320 111454 155668 111486
rect 155320 111218 155376 111454
rect 155612 111218 155668 111454
rect 155320 111134 155668 111218
rect 155320 110898 155376 111134
rect 155612 110898 155668 111134
rect 155320 110866 155668 110898
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 20272 79174 20620 79206
rect 20272 78938 20328 79174
rect 20564 78938 20620 79174
rect 20272 78854 20620 78938
rect 20272 78618 20328 78854
rect 20564 78618 20620 78854
rect 20272 78586 20620 78618
rect 156000 79174 156348 79206
rect 156000 78938 156056 79174
rect 156292 78938 156348 79174
rect 156000 78854 156348 78938
rect 156000 78618 156056 78854
rect 156292 78618 156348 78854
rect 156000 78586 156348 78618
rect 20952 75454 21300 75486
rect 20952 75218 21008 75454
rect 21244 75218 21300 75454
rect 20952 75134 21300 75218
rect 20952 74898 21008 75134
rect 21244 74898 21300 75134
rect 20952 74866 21300 74898
rect 155320 75454 155668 75486
rect 155320 75218 155376 75454
rect 155612 75218 155668 75454
rect 155320 75134 155668 75218
rect 155320 74898 155376 75134
rect 155612 74898 155668 75134
rect 155320 74866 155668 74898
rect 19195 58036 19261 58037
rect 19195 57972 19196 58036
rect 19260 57972 19261 58036
rect 19195 57971 19261 57972
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 36056 50010 36116 50106
rect 37144 50010 37204 50106
rect 35942 49950 36116 50010
rect 37046 49950 37204 50010
rect 38232 50010 38292 50106
rect 39592 50010 39652 50106
rect 40544 50010 40604 50106
rect 38232 49950 38578 50010
rect 39592 49950 39682 50010
rect 18643 47700 18709 47701
rect 18643 47636 18644 47700
rect 18708 47636 18709 47700
rect 18643 47635 18709 47636
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 22054 21014 48064
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 48064
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 48064
rect 35942 47565 36002 49950
rect 37046 48245 37106 49950
rect 37043 48244 37109 48245
rect 37043 48180 37044 48244
rect 37108 48180 37109 48244
rect 37043 48179 37109 48180
rect 35939 47564 36005 47565
rect 35939 47500 35940 47564
rect 36004 47500 36005 47564
rect 35939 47499 36005 47500
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 39454 38414 47940
rect 38518 47837 38578 49950
rect 39622 47973 39682 49950
rect 40542 49950 40604 50010
rect 41768 50010 41828 50106
rect 43128 50010 43188 50106
rect 41768 49950 41890 50010
rect 40542 48109 40602 49950
rect 41830 48109 41890 49950
rect 43118 49950 43188 50010
rect 44216 50010 44276 50106
rect 45440 50010 45500 50106
rect 44216 49950 44282 50010
rect 43118 48245 43178 49950
rect 44222 48245 44282 49950
rect 45326 49950 45500 50010
rect 46528 50010 46588 50106
rect 47616 50010 47676 50106
rect 46528 49950 46674 50010
rect 45326 48245 45386 49950
rect 46614 48245 46674 49950
rect 47534 49950 47676 50010
rect 47534 48245 47594 49950
rect 48296 49605 48356 50106
rect 48704 50010 48764 50106
rect 48638 49950 48764 50010
rect 50064 50010 50124 50106
rect 50064 49950 50170 50010
rect 48293 49604 48359 49605
rect 48293 49540 48294 49604
rect 48358 49540 48359 49604
rect 48293 49539 48359 49540
rect 48638 48245 48698 49950
rect 50110 48245 50170 49950
rect 50744 49605 50804 50106
rect 51288 50010 51348 50106
rect 52376 50010 52436 50106
rect 51288 49950 51458 50010
rect 50741 49604 50807 49605
rect 50741 49540 50742 49604
rect 50806 49540 50807 49604
rect 50741 49539 50807 49540
rect 51398 48245 51458 49950
rect 52318 49950 52436 50010
rect 52318 48245 52378 49950
rect 53464 49877 53524 50106
rect 53461 49876 53527 49877
rect 53461 49812 53462 49876
rect 53526 49812 53527 49876
rect 53461 49811 53527 49812
rect 53600 49605 53660 50106
rect 54552 50010 54612 50106
rect 55912 50010 55972 50106
rect 54526 49950 54612 50010
rect 55814 49950 55972 50010
rect 53597 49604 53663 49605
rect 53597 49540 53598 49604
rect 53662 49540 53663 49604
rect 53597 49539 53663 49540
rect 54526 48245 54586 49950
rect 55814 48245 55874 49950
rect 56048 49605 56108 50106
rect 57000 50010 57060 50106
rect 58088 50010 58148 50106
rect 57000 49950 57162 50010
rect 56045 49604 56111 49605
rect 56045 49540 56046 49604
rect 56110 49540 56111 49604
rect 56045 49539 56111 49540
rect 43115 48244 43181 48245
rect 43115 48180 43116 48244
rect 43180 48180 43181 48244
rect 43115 48179 43181 48180
rect 44219 48244 44285 48245
rect 44219 48180 44220 48244
rect 44284 48180 44285 48244
rect 44219 48179 44285 48180
rect 45323 48244 45389 48245
rect 45323 48180 45324 48244
rect 45388 48180 45389 48244
rect 45323 48179 45389 48180
rect 46611 48244 46677 48245
rect 46611 48180 46612 48244
rect 46676 48180 46677 48244
rect 46611 48179 46677 48180
rect 47531 48244 47597 48245
rect 47531 48180 47532 48244
rect 47596 48180 47597 48244
rect 47531 48179 47597 48180
rect 48635 48244 48701 48245
rect 48635 48180 48636 48244
rect 48700 48180 48701 48244
rect 48635 48179 48701 48180
rect 50107 48244 50173 48245
rect 50107 48180 50108 48244
rect 50172 48180 50173 48244
rect 50107 48179 50173 48180
rect 51395 48244 51461 48245
rect 51395 48180 51396 48244
rect 51460 48180 51461 48244
rect 51395 48179 51461 48180
rect 52315 48244 52381 48245
rect 52315 48180 52316 48244
rect 52380 48180 52381 48244
rect 52315 48179 52381 48180
rect 54523 48244 54589 48245
rect 54523 48180 54524 48244
rect 54588 48180 54589 48244
rect 54523 48179 54589 48180
rect 55811 48244 55877 48245
rect 55811 48180 55812 48244
rect 55876 48180 55877 48244
rect 55811 48179 55877 48180
rect 40539 48108 40605 48109
rect 40539 48044 40540 48108
rect 40604 48044 40605 48108
rect 40539 48043 40605 48044
rect 41827 48108 41893 48109
rect 41827 48044 41828 48108
rect 41892 48044 41893 48108
rect 41827 48043 41893 48044
rect 39619 47972 39685 47973
rect 39619 47908 39620 47972
rect 39684 47908 39685 47972
rect 39619 47907 39685 47908
rect 38515 47836 38581 47837
rect 38515 47772 38516 47836
rect 38580 47772 38581 47836
rect 38515 47771 38581 47772
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 47940
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 46894 45854 47940
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 48064
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 48064
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 47940
rect 57102 47565 57162 49950
rect 58022 49950 58148 50010
rect 58022 48245 58082 49950
rect 58496 49605 58556 50106
rect 59448 50010 59508 50106
rect 59448 49950 59554 50010
rect 58493 49604 58559 49605
rect 58493 49540 58494 49604
rect 58558 49540 58559 49604
rect 58493 49539 58559 49540
rect 59494 48245 59554 49950
rect 60672 49877 60732 50106
rect 61080 50010 61140 50106
rect 61760 50010 61820 50106
rect 62848 50010 62908 50106
rect 61080 49950 61210 50010
rect 60669 49876 60735 49877
rect 60669 49812 60670 49876
rect 60734 49812 60735 49876
rect 60669 49811 60735 49812
rect 61150 48245 61210 49950
rect 61702 49950 61820 50010
rect 62806 49950 62908 50010
rect 63528 50010 63588 50106
rect 63936 50010 63996 50106
rect 65296 50010 65356 50106
rect 65976 50010 66036 50106
rect 66384 50010 66444 50106
rect 67608 50010 67668 50106
rect 63528 49950 63602 50010
rect 61702 48245 61762 49950
rect 62806 48245 62866 49950
rect 63542 48245 63602 49950
rect 63910 49950 63996 50010
rect 65198 49950 65356 50010
rect 65934 49950 66036 50010
rect 66302 49950 66444 50010
rect 67590 49950 67668 50010
rect 68288 50010 68348 50106
rect 68696 50010 68756 50106
rect 68288 49950 68386 50010
rect 58019 48244 58085 48245
rect 58019 48180 58020 48244
rect 58084 48180 58085 48244
rect 58019 48179 58085 48180
rect 59491 48244 59557 48245
rect 59491 48180 59492 48244
rect 59556 48180 59557 48244
rect 59491 48179 59557 48180
rect 61147 48244 61213 48245
rect 61147 48180 61148 48244
rect 61212 48180 61213 48244
rect 61147 48179 61213 48180
rect 61699 48244 61765 48245
rect 61699 48180 61700 48244
rect 61764 48180 61765 48244
rect 61699 48179 61765 48180
rect 62803 48244 62869 48245
rect 62803 48180 62804 48244
rect 62868 48180 62869 48244
rect 62803 48179 62869 48180
rect 63539 48244 63605 48245
rect 63539 48180 63540 48244
rect 63604 48180 63605 48244
rect 63539 48179 63605 48180
rect 63910 48109 63970 49950
rect 65198 48245 65258 49950
rect 65934 48245 65994 49950
rect 66302 48245 66362 49950
rect 67590 48245 67650 49950
rect 68326 48245 68386 49950
rect 68694 49950 68756 50010
rect 69784 50010 69844 50106
rect 71008 50010 71068 50106
rect 69784 49950 69858 50010
rect 68694 48245 68754 49950
rect 69798 48245 69858 49950
rect 70902 49950 71068 50010
rect 70902 48245 70962 49950
rect 71144 49330 71204 50106
rect 72232 50010 72292 50106
rect 73320 50010 73380 50106
rect 71086 49270 71204 49330
rect 72190 49950 72292 50010
rect 73294 49950 73380 50010
rect 73592 50010 73652 50106
rect 74408 50010 74468 50106
rect 73592 49950 73722 50010
rect 65195 48244 65261 48245
rect 65195 48180 65196 48244
rect 65260 48180 65261 48244
rect 65195 48179 65261 48180
rect 65931 48244 65997 48245
rect 65931 48180 65932 48244
rect 65996 48180 65997 48244
rect 65931 48179 65997 48180
rect 66299 48244 66365 48245
rect 66299 48180 66300 48244
rect 66364 48180 66365 48244
rect 66299 48179 66365 48180
rect 67587 48244 67653 48245
rect 67587 48180 67588 48244
rect 67652 48180 67653 48244
rect 67587 48179 67653 48180
rect 68323 48244 68389 48245
rect 68323 48180 68324 48244
rect 68388 48180 68389 48244
rect 68323 48179 68389 48180
rect 68691 48244 68757 48245
rect 68691 48180 68692 48244
rect 68756 48180 68757 48244
rect 68691 48179 68757 48180
rect 69795 48244 69861 48245
rect 69795 48180 69796 48244
rect 69860 48180 69861 48244
rect 69795 48179 69861 48180
rect 70899 48244 70965 48245
rect 70899 48180 70900 48244
rect 70964 48180 70965 48244
rect 70899 48179 70965 48180
rect 71086 48109 71146 49270
rect 72190 48245 72250 49950
rect 73294 48245 73354 49950
rect 73662 48245 73722 49950
rect 74398 49950 74468 50010
rect 74398 48245 74458 49950
rect 75768 49710 75828 50106
rect 75686 49650 75828 49710
rect 76040 49710 76100 50106
rect 76992 49710 77052 50106
rect 78080 49710 78140 50106
rect 78488 49710 78548 50106
rect 76040 49650 76114 49710
rect 72187 48244 72253 48245
rect 72187 48180 72188 48244
rect 72252 48180 72253 48244
rect 72187 48179 72253 48180
rect 73291 48244 73357 48245
rect 73291 48180 73292 48244
rect 73356 48180 73357 48244
rect 73291 48179 73357 48180
rect 73659 48244 73725 48245
rect 73659 48180 73660 48244
rect 73724 48180 73725 48244
rect 73659 48179 73725 48180
rect 74395 48244 74461 48245
rect 74395 48180 74396 48244
rect 74460 48180 74461 48244
rect 74395 48179 74461 48180
rect 63907 48108 63973 48109
rect 63907 48044 63908 48108
rect 63972 48044 63973 48108
rect 63907 48043 63973 48044
rect 71083 48108 71149 48109
rect 71083 48044 71084 48108
rect 71148 48044 71149 48108
rect 71083 48043 71149 48044
rect 57099 47564 57165 47565
rect 57099 47500 57100 47564
rect 57164 47500 57165 47564
rect 57099 47499 57165 47500
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 47940
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 29494 64454 47940
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 47940
rect 75686 47565 75746 49650
rect 76054 48245 76114 49650
rect 76974 49650 77052 49710
rect 78078 49650 78140 49710
rect 78446 49650 78548 49710
rect 79168 49710 79228 50106
rect 79168 49650 79242 49710
rect 76974 48245 77034 49650
rect 78078 48245 78138 49650
rect 78446 48245 78506 49650
rect 76051 48244 76117 48245
rect 76051 48180 76052 48244
rect 76116 48180 76117 48244
rect 76051 48179 76117 48180
rect 76971 48244 77037 48245
rect 76971 48180 76972 48244
rect 77036 48180 77037 48244
rect 76971 48179 77037 48180
rect 78075 48244 78141 48245
rect 78075 48180 78076 48244
rect 78140 48180 78141 48244
rect 78075 48179 78141 48180
rect 78443 48244 78509 48245
rect 78443 48180 78444 48244
rect 78508 48180 78509 48244
rect 78443 48179 78509 48180
rect 79182 47973 79242 49650
rect 80936 49605 80996 50106
rect 83520 49605 83580 50106
rect 85968 49605 86028 50106
rect 88280 49605 88340 50106
rect 91000 49741 91060 50106
rect 93448 50010 93508 50106
rect 93448 49950 93594 50010
rect 90997 49740 91063 49741
rect 90997 49676 90998 49740
rect 91062 49676 91063 49740
rect 90997 49675 91063 49676
rect 80933 49604 80999 49605
rect 80933 49540 80934 49604
rect 80998 49540 80999 49604
rect 80933 49539 80999 49540
rect 83517 49604 83583 49605
rect 83517 49540 83518 49604
rect 83582 49540 83583 49604
rect 83517 49539 83583 49540
rect 85965 49604 86031 49605
rect 85965 49540 85966 49604
rect 86030 49540 86031 49604
rect 85965 49539 86031 49540
rect 88277 49604 88343 49605
rect 88277 49540 88278 49604
rect 88342 49540 88343 49604
rect 88277 49539 88343 49540
rect 93534 48245 93594 49950
rect 95896 49741 95956 50106
rect 95893 49740 95959 49741
rect 95893 49676 95894 49740
rect 95958 49676 95959 49740
rect 95893 49675 95959 49676
rect 98480 49605 98540 50106
rect 100928 50010 100988 50106
rect 100894 49950 100988 50010
rect 98477 49604 98543 49605
rect 98477 49540 98478 49604
rect 98542 49540 98543 49604
rect 98477 49539 98543 49540
rect 100894 48245 100954 49950
rect 103512 49605 103572 50106
rect 105960 49605 106020 50106
rect 108544 50010 108604 50106
rect 110992 50010 111052 50106
rect 113440 50010 113500 50106
rect 115888 50010 115948 50106
rect 108544 49950 108682 50010
rect 110992 49950 111074 50010
rect 103509 49604 103575 49605
rect 103509 49540 103510 49604
rect 103574 49540 103575 49604
rect 103509 49539 103575 49540
rect 105957 49604 106023 49605
rect 105957 49540 105958 49604
rect 106022 49540 106023 49604
rect 105957 49539 106023 49540
rect 108622 48245 108682 49950
rect 111014 48245 111074 49950
rect 113406 49950 113500 50010
rect 115798 49950 115948 50010
rect 118472 50010 118532 50106
rect 118472 49950 118618 50010
rect 113406 49469 113466 49950
rect 113403 49468 113469 49469
rect 113403 49404 113404 49468
rect 113468 49404 113469 49468
rect 113403 49403 113469 49404
rect 115798 48245 115858 49950
rect 118558 48245 118618 49950
rect 120920 49605 120980 50106
rect 123368 50010 123428 50106
rect 125952 50010 126012 50106
rect 123342 49950 123428 50010
rect 125918 49950 126012 50010
rect 120917 49604 120983 49605
rect 120917 49540 120918 49604
rect 120982 49540 120983 49604
rect 120917 49539 120983 49540
rect 93531 48244 93597 48245
rect 93531 48180 93532 48244
rect 93596 48180 93597 48244
rect 93531 48179 93597 48180
rect 100891 48244 100957 48245
rect 100891 48180 100892 48244
rect 100956 48180 100957 48244
rect 100891 48179 100957 48180
rect 108619 48244 108685 48245
rect 108619 48180 108620 48244
rect 108684 48180 108685 48244
rect 108619 48179 108685 48180
rect 111011 48244 111077 48245
rect 111011 48180 111012 48244
rect 111076 48180 111077 48244
rect 111011 48179 111077 48180
rect 115795 48244 115861 48245
rect 115795 48180 115796 48244
rect 115860 48180 115861 48244
rect 115795 48179 115861 48180
rect 118555 48244 118621 48245
rect 118555 48180 118556 48244
rect 118620 48180 118621 48244
rect 118555 48179 118621 48180
rect 123342 48109 123402 49950
rect 125918 48245 125978 49950
rect 125915 48244 125981 48245
rect 125915 48180 125916 48244
rect 125980 48180 125981 48244
rect 125915 48179 125981 48180
rect 123339 48108 123405 48109
rect 79179 47972 79245 47973
rect 75683 47564 75749 47565
rect 75683 47500 75684 47564
rect 75748 47500 75749 47564
rect 75683 47499 75749 47500
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 47940
rect 79179 47908 79180 47972
rect 79244 47908 79245 47972
rect 79179 47907 79245 47908
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 48064
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 48064
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 48064
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 48064
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 48064
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 48064
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 48064
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 47940
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 48064
rect 123339 48044 123340 48108
rect 123404 48044 123405 48108
rect 123339 48043 123405 48044
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 47940
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 48064
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 48064
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 48064
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 48064
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 48064
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 48064
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 48064
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 48064
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 490054 165014 525498
rect 164394 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 165014 490054
rect 164394 489734 165014 489818
rect 164394 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 165014 489734
rect 164394 454054 165014 489498
rect 164394 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 165014 454054
rect 164394 453734 165014 453818
rect 164394 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 165014 453734
rect 164394 418054 165014 453498
rect 164394 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 165014 418054
rect 164394 417734 165014 417818
rect 164394 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 165014 417734
rect 164394 382054 165014 417498
rect 164394 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 165014 382054
rect 164394 381734 165014 381818
rect 164394 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 165014 381734
rect 164394 346054 165014 381498
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 168114 601774 168734 637218
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 168114 565774 168734 601218
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 168114 529774 168734 565218
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 168114 493774 168734 529218
rect 168114 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 168734 493774
rect 168114 493454 168734 493538
rect 168114 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 168734 493454
rect 168114 457774 168734 493218
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 168114 421774 168734 457218
rect 168114 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 168734 421774
rect 168114 421454 168734 421538
rect 168114 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 168734 421454
rect 168114 385774 168734 421218
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 168114 349774 168734 385218
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 168114 241774 168734 277218
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 168114 61774 168734 97218
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 168114 25774 168734 61218
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 171834 569494 172454 604938
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 171834 533494 172454 568938
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 171834 497494 172454 532938
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 171834 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 172454 497494
rect 171834 497174 172454 497258
rect 171834 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 172454 497174
rect 171834 461494 172454 496938
rect 171834 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 172454 461494
rect 171834 461174 172454 461258
rect 171834 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 172454 461174
rect 171834 425494 172454 460938
rect 171834 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 172454 425494
rect 171834 425174 172454 425258
rect 171834 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 172454 425174
rect 171834 389494 172454 424938
rect 171834 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 172454 389494
rect 171834 389174 172454 389258
rect 171834 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 172454 389174
rect 171834 353494 172454 388938
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 171834 245494 172454 280938
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 171834 101494 172454 136938
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 171834 65494 172454 100938
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 186267 682004 186333 682005
rect 186267 681940 186268 682004
rect 186332 681940 186333 682004
rect 186267 681939 186333 681940
rect 186270 678197 186330 681939
rect 186267 678196 186333 678197
rect 186267 678132 186268 678196
rect 186332 678132 186333 678196
rect 186267 678131 186333 678132
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 658894 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 679452 193574 698058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 193811 682140 193877 682141
rect 193811 682076 193812 682140
rect 193876 682076 193877 682140
rect 193811 682075 193877 682076
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 192954 482614 193574 500068
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192339 453116 192405 453117
rect 192339 453052 192340 453116
rect 192404 453052 192405 453116
rect 192339 453051 192405 453052
rect 191603 452708 191669 452709
rect 191603 452644 191604 452708
rect 191668 452644 191669 452708
rect 191603 452643 191669 452644
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 191606 250477 191666 452643
rect 192342 347173 192402 453051
rect 192954 446614 193574 482058
rect 193814 457469 193874 682075
rect 193995 681868 194061 681869
rect 193995 681804 193996 681868
rect 194060 681804 194061 681868
rect 193995 681803 194061 681804
rect 193998 462909 194058 681803
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 196674 594334 197294 629778
rect 196674 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 197294 594334
rect 196674 594014 197294 594098
rect 196674 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 197294 594014
rect 196674 558334 197294 593778
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 196674 486334 197294 521778
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 193995 462908 194061 462909
rect 193995 462844 193996 462908
rect 194060 462844 194061 462908
rect 193995 462843 194061 462844
rect 193811 457468 193877 457469
rect 193811 457404 193812 457468
rect 193876 457404 193877 457468
rect 193811 457403 193877 457404
rect 193995 450396 194061 450397
rect 193995 450332 193996 450396
rect 194060 450332 194061 450396
rect 193995 450331 194061 450332
rect 196674 450334 197294 485778
rect 193811 449308 193877 449309
rect 193811 449244 193812 449308
rect 193876 449244 193877 449308
rect 193811 449243 193877 449244
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192339 347172 192405 347173
rect 192339 347108 192340 347172
rect 192404 347108 192405 347172
rect 192339 347107 192405 347108
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 191603 250476 191669 250477
rect 191603 250412 191604 250476
rect 191668 250412 191669 250476
rect 191603 250411 191669 250412
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 193814 31789 193874 449243
rect 193811 31788 193877 31789
rect 193811 31724 193812 31788
rect 193876 31724 193877 31788
rect 193811 31723 193877 31724
rect 193998 19413 194058 450331
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 194208 435454 194528 435486
rect 194208 435218 194250 435454
rect 194486 435218 194528 435454
rect 194208 435134 194528 435218
rect 194208 434898 194250 435134
rect 194486 434898 194528 435134
rect 194208 434866 194528 434898
rect 196674 414334 197294 449778
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 194208 399454 194528 399486
rect 194208 399218 194250 399454
rect 194486 399218 194528 399454
rect 194208 399134 194528 399218
rect 194208 398898 194250 399134
rect 194486 398898 194528 399134
rect 194208 398866 194528 398898
rect 196674 378334 197294 413778
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 194208 363454 194528 363486
rect 194208 363218 194250 363454
rect 194486 363218 194528 363454
rect 194208 363134 194528 363218
rect 194208 362898 194250 363134
rect 194486 362898 194528 363134
rect 194208 362866 194528 362898
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 194208 327454 194528 327486
rect 194208 327218 194250 327454
rect 194486 327218 194528 327454
rect 194208 327134 194528 327218
rect 194208 326898 194250 327134
rect 194486 326898 194528 327134
rect 194208 326866 194528 326898
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 194208 291454 194528 291486
rect 194208 291218 194250 291454
rect 194486 291218 194528 291454
rect 194208 291134 194528 291218
rect 194208 290898 194250 291134
rect 194486 290898 194528 291134
rect 194208 290866 194528 290898
rect 196674 270334 197294 305778
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 194208 255454 194528 255486
rect 194208 255218 194250 255454
rect 194486 255218 194528 255454
rect 194208 255134 194528 255218
rect 194208 254898 194250 255134
rect 194486 254898 194528 255134
rect 194208 254866 194528 254898
rect 196674 234334 197294 269778
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 198334 197294 233778
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 196674 162334 197294 197778
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 196674 90334 197294 125778
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 196674 54334 197294 89778
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 193995 19412 194061 19413
rect 193995 19348 193996 19412
rect 194060 19348 194061 19412
rect 193995 19347 194061 19348
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 598054 201014 633498
rect 200394 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 201014 598054
rect 200394 597734 201014 597818
rect 200394 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 201014 597734
rect 200394 562054 201014 597498
rect 200394 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 201014 562054
rect 200394 561734 201014 561818
rect 200394 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 201014 561734
rect 200394 526054 201014 561498
rect 200394 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 201014 526054
rect 200394 525734 201014 525818
rect 200394 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 201014 525734
rect 200394 490054 201014 525498
rect 200394 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 201014 490054
rect 200394 489734 201014 489818
rect 200394 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 201014 489734
rect 200394 454054 201014 489498
rect 200394 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 201014 454054
rect 200394 453734 201014 453818
rect 200394 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 201014 453734
rect 200394 418054 201014 453498
rect 200394 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 201014 418054
rect 200394 417734 201014 417818
rect 200394 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 201014 417734
rect 200394 382054 201014 417498
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 274054 201014 309498
rect 200394 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 201014 274054
rect 200394 273734 201014 273818
rect 200394 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 201014 273734
rect 200394 238054 201014 273498
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 202054 201014 237498
rect 200394 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 201014 202054
rect 200394 201734 201014 201818
rect 200394 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 201014 201734
rect 200394 166054 201014 201498
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 200394 94054 201014 129498
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 200394 58054 201014 93498
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 601774 204734 637218
rect 204114 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 204734 601774
rect 204114 601454 204734 601538
rect 204114 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 204734 601454
rect 204114 565774 204734 601218
rect 204114 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 204734 565774
rect 204114 565454 204734 565538
rect 204114 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 204734 565454
rect 204114 529774 204734 565218
rect 204114 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 204734 529774
rect 204114 529454 204734 529538
rect 204114 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 204734 529454
rect 204114 493774 204734 529218
rect 204114 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 204734 493774
rect 204114 493454 204734 493538
rect 204114 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 204734 493454
rect 204114 457774 204734 493218
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 204114 421774 204734 457218
rect 204114 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 204734 421774
rect 204114 421454 204734 421538
rect 204114 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 204734 421454
rect 204114 385774 204734 421218
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 204114 277774 204734 313218
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 204114 241774 204734 277218
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 205774 204734 241218
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 204114 169774 204734 205218
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 204114 97774 204734 133218
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 204114 61774 204734 97218
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 605494 208454 640938
rect 207834 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 208454 605494
rect 207834 605174 208454 605258
rect 207834 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 208454 605174
rect 207834 569494 208454 604938
rect 207834 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 208454 569494
rect 207834 569174 208454 569258
rect 207834 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 208454 569174
rect 207834 533494 208454 568938
rect 207834 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 208454 533494
rect 207834 533174 208454 533258
rect 207834 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 208454 533174
rect 207834 497494 208454 532938
rect 207834 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 208454 497494
rect 207834 497174 208454 497258
rect 207834 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 208454 497174
rect 207834 461494 208454 496938
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 207834 425494 208454 460938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 209568 439174 209888 439206
rect 209568 438938 209610 439174
rect 209846 438938 209888 439174
rect 209568 438854 209888 438938
rect 209568 438618 209610 438854
rect 209846 438618 209888 438854
rect 209568 438586 209888 438618
rect 207834 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 208454 425494
rect 207834 425174 208454 425258
rect 207834 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 208454 425174
rect 207834 389494 208454 424938
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 209568 403174 209888 403206
rect 209568 402938 209610 403174
rect 209846 402938 209888 403174
rect 209568 402854 209888 402938
rect 209568 402618 209610 402854
rect 209846 402618 209888 402854
rect 209568 402586 209888 402618
rect 207834 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 208454 389494
rect 207834 389174 208454 389258
rect 207834 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 208454 389174
rect 207834 353494 208454 388938
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 209568 367174 209888 367206
rect 209568 366938 209610 367174
rect 209846 366938 209888 367174
rect 209568 366854 209888 366938
rect 209568 366618 209610 366854
rect 209846 366618 209888 366854
rect 209568 366586 209888 366618
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 209568 331174 209888 331206
rect 209568 330938 209610 331174
rect 209846 330938 209888 331174
rect 209568 330854 209888 330938
rect 209568 330618 209610 330854
rect 209846 330618 209888 330854
rect 209568 330586 209888 330618
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 207834 281494 208454 316938
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 209568 295174 209888 295206
rect 209568 294938 209610 295174
rect 209846 294938 209888 295174
rect 209568 294854 209888 294938
rect 209568 294618 209610 294854
rect 209846 294618 209888 294854
rect 209568 294586 209888 294618
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 207834 245494 208454 280938
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 209568 259174 209888 259206
rect 209568 258938 209610 259174
rect 209846 258938 209888 259174
rect 209568 258854 209888 258938
rect 209568 258618 209610 258854
rect 209846 258618 209888 258854
rect 209568 258586 209888 258618
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 209494 208454 244938
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 207834 173494 208454 208938
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 101494 208454 136938
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 207834 65494 208454 100938
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 449580 225854 478338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 224928 435454 225248 435486
rect 224928 435218 224970 435454
rect 225206 435218 225248 435454
rect 224928 435134 225248 435218
rect 224928 434898 224970 435134
rect 225206 434898 225248 435134
rect 224928 434866 225248 434898
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 224928 399454 225248 399486
rect 224928 399218 224970 399454
rect 225206 399218 225248 399454
rect 224928 399134 225248 399218
rect 224928 398898 224970 399134
rect 225206 398898 225248 399134
rect 224928 398866 225248 398898
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 224928 363454 225248 363486
rect 224928 363218 224970 363454
rect 225206 363218 225248 363454
rect 224928 363134 225248 363218
rect 224928 362898 224970 363134
rect 225206 362898 225248 363134
rect 224928 362866 225248 362898
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 224928 327454 225248 327486
rect 224928 327218 224970 327454
rect 225206 327218 225248 327454
rect 224928 327134 225248 327218
rect 224928 326898 224970 327134
rect 225206 326898 225248 327134
rect 224928 326866 225248 326898
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 224928 291454 225248 291486
rect 224928 291218 224970 291454
rect 225206 291218 225248 291454
rect 224928 291134 225248 291218
rect 224928 290898 224970 291134
rect 225206 290898 225248 291134
rect 224928 290866 225248 290898
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 224928 255454 225248 255486
rect 224928 255218 224970 255454
rect 225206 255218 225248 255454
rect 224928 255134 225248 255218
rect 224928 254898 224970 255134
rect 225206 254898 225248 255134
rect 224928 254866 225248 254898
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 226894 225854 250068
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 630334 233294 665778
rect 232674 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 233294 630334
rect 232674 630014 233294 630098
rect 232674 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 233294 630014
rect 232674 594334 233294 629778
rect 232674 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 233294 594334
rect 232674 594014 233294 594098
rect 232674 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 233294 594014
rect 232674 558334 233294 593778
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 232674 522334 233294 557778
rect 232674 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 233294 522334
rect 232674 522014 233294 522098
rect 232674 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 233294 522014
rect 232674 486334 233294 521778
rect 232674 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 233294 486334
rect 232674 486014 233294 486098
rect 232674 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 233294 486014
rect 232674 450334 233294 485778
rect 232674 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 233294 450334
rect 232674 450014 233294 450098
rect 232674 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 233294 450014
rect 232674 414334 233294 449778
rect 232674 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 233294 414334
rect 232674 414014 233294 414098
rect 232674 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 233294 414014
rect 232674 378334 233294 413778
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 232674 342334 233294 377778
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232674 306334 233294 341778
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232674 270334 233294 305778
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 232674 234334 233294 269778
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 232674 198334 233294 233778
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 232674 162334 233294 197778
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232674 126334 233294 161778
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 90334 233294 125778
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 232674 54334 233294 89778
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 598054 237014 633498
rect 236394 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 237014 598054
rect 236394 597734 237014 597818
rect 236394 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 237014 597734
rect 236394 562054 237014 597498
rect 236394 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 237014 562054
rect 236394 561734 237014 561818
rect 236394 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 237014 561734
rect 236394 526054 237014 561498
rect 236394 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 237014 526054
rect 236394 525734 237014 525818
rect 236394 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 237014 525734
rect 236394 490054 237014 525498
rect 236394 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 237014 490054
rect 236394 489734 237014 489818
rect 236394 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 237014 489734
rect 236394 454054 237014 489498
rect 236394 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 237014 454054
rect 236394 453734 237014 453818
rect 236394 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 237014 453734
rect 236394 418054 237014 453498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 601774 240734 637218
rect 240114 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 240734 601774
rect 240114 601454 240734 601538
rect 240114 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 240734 601454
rect 240114 565774 240734 601218
rect 240114 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 240734 565774
rect 240114 565454 240734 565538
rect 240114 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 240734 565454
rect 240114 529774 240734 565218
rect 240114 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 240734 529774
rect 240114 529454 240734 529538
rect 240114 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 240734 529454
rect 240114 493774 240734 529218
rect 240114 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 240734 493774
rect 240114 493454 240734 493538
rect 240114 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 240734 493454
rect 240114 457774 240734 493218
rect 240114 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 240734 457774
rect 240114 457454 240734 457538
rect 240114 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 240734 457454
rect 240114 449580 240734 457218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 605494 244454 640938
rect 243834 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 244454 605494
rect 243834 605174 244454 605258
rect 243834 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 244454 605174
rect 243834 569494 244454 604938
rect 243834 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 244454 569494
rect 243834 569174 244454 569258
rect 243834 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 244454 569174
rect 243834 533494 244454 568938
rect 243834 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 244454 533494
rect 243834 533174 244454 533258
rect 243834 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 244454 533174
rect 243834 497494 244454 532938
rect 243834 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 244454 497494
rect 243834 497174 244454 497258
rect 243834 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 244454 497174
rect 243834 461494 244454 496938
rect 243834 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 244454 461494
rect 243834 461174 244454 461258
rect 243834 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 244454 461174
rect 240288 439174 240608 439206
rect 240288 438938 240330 439174
rect 240566 438938 240608 439174
rect 240288 438854 240608 438938
rect 240288 438618 240330 438854
rect 240566 438618 240608 438854
rect 240288 438586 240608 438618
rect 236394 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 237014 418054
rect 236394 417734 237014 417818
rect 236394 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 237014 417734
rect 236394 382054 237014 417498
rect 243834 425494 244454 460938
rect 243834 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 244454 425494
rect 243834 425174 244454 425258
rect 243834 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 244454 425174
rect 240288 403174 240608 403206
rect 240288 402938 240330 403174
rect 240566 402938 240608 403174
rect 240288 402854 240608 402938
rect 240288 402618 240330 402854
rect 240566 402618 240608 402854
rect 240288 402586 240608 402618
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 236394 346054 237014 381498
rect 243834 389494 244454 424938
rect 243834 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 244454 389494
rect 243834 389174 244454 389258
rect 243834 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 244454 389174
rect 240288 367174 240608 367206
rect 240288 366938 240330 367174
rect 240566 366938 240608 367174
rect 240288 366854 240608 366938
rect 240288 366618 240330 366854
rect 240566 366618 240608 366854
rect 240288 366586 240608 366618
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 236394 310054 237014 345498
rect 243834 353494 244454 388938
rect 243834 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 244454 353494
rect 243834 353174 244454 353258
rect 243834 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 244454 353174
rect 240288 331174 240608 331206
rect 240288 330938 240330 331174
rect 240566 330938 240608 331174
rect 240288 330854 240608 330938
rect 240288 330618 240330 330854
rect 240566 330618 240608 330854
rect 240288 330586 240608 330618
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 236394 274054 237014 309498
rect 243834 317494 244454 352938
rect 243834 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 244454 317494
rect 243834 317174 244454 317258
rect 243834 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 244454 317174
rect 240288 295174 240608 295206
rect 240288 294938 240330 295174
rect 240566 294938 240608 295174
rect 240288 294854 240608 294938
rect 240288 294618 240330 294854
rect 240566 294618 240608 294854
rect 240288 294586 240608 294618
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 236394 238054 237014 273498
rect 243834 281494 244454 316938
rect 243834 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 244454 281494
rect 243834 281174 244454 281258
rect 243834 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 244454 281174
rect 240288 259174 240608 259206
rect 240288 258938 240330 259174
rect 240566 258938 240608 259174
rect 240288 258854 240608 258938
rect 240288 258618 240330 258854
rect 240566 258618 240608 258854
rect 240288 258586 240608 258618
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 236394 202054 237014 237498
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 236394 166054 237014 201498
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 236394 130054 237014 165498
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 236394 94054 237014 129498
rect 236394 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 237014 94054
rect 236394 93734 237014 93818
rect 236394 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 237014 93734
rect 236394 58054 237014 93498
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 241774 240734 250068
rect 240114 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 240734 241774
rect 240114 241454 240734 241538
rect 240114 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 240734 241454
rect 240114 205774 240734 241218
rect 240114 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 240734 205774
rect 240114 205454 240734 205538
rect 240114 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 240734 205454
rect 240114 169774 240734 205218
rect 240114 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 240734 169774
rect 240114 169454 240734 169538
rect 240114 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 240734 169454
rect 240114 133774 240734 169218
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 240114 97774 240734 133218
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 240114 61774 240734 97218
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 245494 244454 280938
rect 243834 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 244454 245494
rect 243834 245174 244454 245258
rect 243834 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 244454 245174
rect 243834 209494 244454 244938
rect 243834 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 244454 209494
rect 243834 209174 244454 209258
rect 243834 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 244454 209174
rect 243834 173494 244454 208938
rect 243834 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 244454 173494
rect 243834 173174 244454 173258
rect 243834 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 244454 173174
rect 243834 137494 244454 172938
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 243834 101494 244454 136938
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 243834 65494 244454 100938
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 451537 258134 474618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 451537 261854 478338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 451537 265574 482058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 630334 269294 665778
rect 268674 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 269294 630334
rect 268674 630014 269294 630098
rect 268674 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 269294 630014
rect 268674 594334 269294 629778
rect 268674 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 269294 594334
rect 268674 594014 269294 594098
rect 268674 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 269294 594014
rect 268674 558334 269294 593778
rect 268674 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 269294 558334
rect 268674 558014 269294 558098
rect 268674 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 269294 558014
rect 268674 522334 269294 557778
rect 268674 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 269294 522334
rect 268674 522014 269294 522098
rect 268674 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 269294 522014
rect 268674 486334 269294 521778
rect 268674 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 269294 486334
rect 268674 486014 269294 486098
rect 268674 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 269294 486014
rect 268674 451537 269294 485778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 634054 273014 669498
rect 272394 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 273014 634054
rect 272394 633734 273014 633818
rect 272394 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 273014 633734
rect 272394 598054 273014 633498
rect 272394 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 273014 598054
rect 272394 597734 273014 597818
rect 272394 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 273014 597734
rect 272394 562054 273014 597498
rect 272394 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 273014 562054
rect 272394 561734 273014 561818
rect 272394 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 273014 561734
rect 272394 526054 273014 561498
rect 272394 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 273014 526054
rect 272394 525734 273014 525818
rect 272394 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 273014 525734
rect 272394 490054 273014 525498
rect 272394 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 273014 490054
rect 272394 489734 273014 489818
rect 272394 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 273014 489734
rect 272394 454054 273014 489498
rect 272394 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 273014 454054
rect 272394 453734 273014 453818
rect 272394 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 273014 453734
rect 272394 451537 273014 453498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 637774 276734 673218
rect 276114 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 276734 637774
rect 276114 637454 276734 637538
rect 276114 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 276734 637454
rect 276114 601774 276734 637218
rect 276114 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 276734 601774
rect 276114 601454 276734 601538
rect 276114 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 276734 601454
rect 276114 565774 276734 601218
rect 276114 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 276734 565774
rect 276114 565454 276734 565538
rect 276114 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 276734 565454
rect 276114 529774 276734 565218
rect 276114 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 276734 529774
rect 276114 529454 276734 529538
rect 276114 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 276734 529454
rect 276114 493774 276734 529218
rect 276114 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 276734 493774
rect 276114 493454 276734 493538
rect 276114 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 276734 493454
rect 276114 457774 276734 493218
rect 276114 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 276734 457774
rect 276114 457454 276734 457538
rect 276114 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 276734 457454
rect 276114 451537 276734 457218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 641494 280454 676938
rect 279834 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 280454 641494
rect 279834 641174 280454 641258
rect 279834 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 280454 641174
rect 279834 605494 280454 640938
rect 279834 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 280454 605494
rect 279834 605174 280454 605258
rect 279834 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 280454 605174
rect 279834 569494 280454 604938
rect 279834 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 280454 569494
rect 279834 569174 280454 569258
rect 279834 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 280454 569174
rect 279834 533494 280454 568938
rect 279834 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 280454 533494
rect 279834 533174 280454 533258
rect 279834 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 280454 533174
rect 279834 497494 280454 532938
rect 279834 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 280454 497494
rect 279834 497174 280454 497258
rect 279834 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 280454 497174
rect 279834 461494 280454 496938
rect 279834 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 280454 461494
rect 279834 461174 280454 461258
rect 279834 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 280454 461174
rect 279834 451537 280454 460938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 451537 290414 470898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 451537 294134 474618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 451537 297854 478338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 451537 301574 482058
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 630334 305294 665778
rect 304674 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 305294 630334
rect 304674 630014 305294 630098
rect 304674 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 305294 630014
rect 304674 594334 305294 629778
rect 304674 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 305294 594334
rect 304674 594014 305294 594098
rect 304674 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 305294 594014
rect 304674 558334 305294 593778
rect 304674 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 305294 558334
rect 304674 558014 305294 558098
rect 304674 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 305294 558014
rect 304674 522334 305294 557778
rect 304674 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 305294 522334
rect 304674 522014 305294 522098
rect 304674 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 305294 522014
rect 304674 486334 305294 521778
rect 304674 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 305294 486334
rect 304674 486014 305294 486098
rect 304674 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 305294 486014
rect 304674 451537 305294 485778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 634054 309014 669498
rect 308394 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 309014 634054
rect 308394 633734 309014 633818
rect 308394 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 309014 633734
rect 308394 598054 309014 633498
rect 308394 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 309014 598054
rect 308394 597734 309014 597818
rect 308394 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 309014 597734
rect 308394 562054 309014 597498
rect 308394 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 309014 562054
rect 308394 561734 309014 561818
rect 308394 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 309014 561734
rect 308394 526054 309014 561498
rect 308394 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 309014 526054
rect 308394 525734 309014 525818
rect 308394 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 309014 525734
rect 308394 490054 309014 525498
rect 308394 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 309014 490054
rect 308394 489734 309014 489818
rect 308394 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 309014 489734
rect 308394 454054 309014 489498
rect 308394 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 309014 454054
rect 308394 453734 309014 453818
rect 308394 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 309014 453734
rect 308394 451537 309014 453498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 637774 312734 673218
rect 312114 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 312734 637774
rect 312114 637454 312734 637538
rect 312114 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 312734 637454
rect 312114 601774 312734 637218
rect 312114 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 312734 601774
rect 312114 601454 312734 601538
rect 312114 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 312734 601454
rect 312114 565774 312734 601218
rect 312114 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 312734 565774
rect 312114 565454 312734 565538
rect 312114 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 312734 565454
rect 312114 529774 312734 565218
rect 312114 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 312734 529774
rect 312114 529454 312734 529538
rect 312114 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 312734 529454
rect 312114 493774 312734 529218
rect 312114 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 312734 493774
rect 312114 493454 312734 493538
rect 312114 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 312734 493454
rect 312114 457774 312734 493218
rect 312114 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 312734 457774
rect 312114 457454 312734 457538
rect 312114 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 312734 457454
rect 312114 451537 312734 457218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 641494 316454 676938
rect 315834 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 316454 641494
rect 315834 641174 316454 641258
rect 315834 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 316454 641174
rect 315834 605494 316454 640938
rect 315834 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 316454 605494
rect 315834 605174 316454 605258
rect 315834 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 316454 605174
rect 315834 569494 316454 604938
rect 315834 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 316454 569494
rect 315834 569174 316454 569258
rect 315834 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 316454 569174
rect 315834 533494 316454 568938
rect 315834 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 316454 533494
rect 315834 533174 316454 533258
rect 315834 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 316454 533174
rect 315834 497494 316454 532938
rect 315834 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 316454 497494
rect 315834 497174 316454 497258
rect 315834 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 316454 497174
rect 315834 461494 316454 496938
rect 315834 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 316454 461494
rect 315834 461174 316454 461258
rect 315834 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 316454 461174
rect 315834 451537 316454 460938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 451537 326414 470898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 451537 330134 474618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 451537 333854 478338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 451537 337574 482058
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 630334 341294 665778
rect 340674 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 341294 630334
rect 340674 630014 341294 630098
rect 340674 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 341294 630014
rect 340674 594334 341294 629778
rect 340674 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 341294 594334
rect 340674 594014 341294 594098
rect 340674 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 341294 594014
rect 340674 558334 341294 593778
rect 340674 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 341294 558334
rect 340674 558014 341294 558098
rect 340674 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 341294 558014
rect 340674 522334 341294 557778
rect 340674 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 341294 522334
rect 340674 522014 341294 522098
rect 340674 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 341294 522014
rect 340674 486334 341294 521778
rect 340674 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 341294 486334
rect 340674 486014 341294 486098
rect 340674 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 341294 486014
rect 340674 451537 341294 485778
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 344394 598054 345014 633498
rect 344394 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 345014 598054
rect 344394 597734 345014 597818
rect 344394 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 345014 597734
rect 344394 562054 345014 597498
rect 344394 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 345014 562054
rect 344394 561734 345014 561818
rect 344394 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 345014 561734
rect 344394 526054 345014 561498
rect 344394 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 345014 526054
rect 344394 525734 345014 525818
rect 344394 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 345014 525734
rect 344394 490054 345014 525498
rect 344394 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 345014 490054
rect 344394 489734 345014 489818
rect 344394 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 345014 489734
rect 344394 454054 345014 489498
rect 344394 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 345014 454054
rect 344394 453734 345014 453818
rect 344394 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 345014 453734
rect 344394 451537 345014 453498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 601774 348734 637218
rect 348114 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 348734 601774
rect 348114 601454 348734 601538
rect 348114 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 348734 601454
rect 348114 565774 348734 601218
rect 348114 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 348734 565774
rect 348114 565454 348734 565538
rect 348114 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 348734 565454
rect 348114 529774 348734 565218
rect 348114 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 348734 529774
rect 348114 529454 348734 529538
rect 348114 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 348734 529454
rect 348114 493774 348734 529218
rect 348114 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 348734 493774
rect 348114 493454 348734 493538
rect 348114 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 348734 493454
rect 348114 457774 348734 493218
rect 348114 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 348734 457774
rect 348114 457454 348734 457538
rect 348114 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 348734 457454
rect 348114 451537 348734 457218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 605494 352454 640938
rect 351834 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 352454 605494
rect 351834 605174 352454 605258
rect 351834 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 352454 605174
rect 351834 569494 352454 604938
rect 351834 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 352454 569494
rect 351834 569174 352454 569258
rect 351834 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 352454 569174
rect 351834 533494 352454 568938
rect 351834 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 352454 533494
rect 351834 533174 352454 533258
rect 351834 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 352454 533174
rect 351834 497494 352454 532938
rect 351834 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 352454 497494
rect 351834 497174 352454 497258
rect 351834 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 352454 497174
rect 351834 461494 352454 496938
rect 351834 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 352454 461494
rect 351834 461174 352454 461258
rect 351834 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 352454 461174
rect 351834 451537 352454 460938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 451537 362414 470898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 451537 366134 474618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 271008 439174 271328 439206
rect 271008 438938 271050 439174
rect 271286 438938 271328 439174
rect 271008 438854 271328 438938
rect 271008 438618 271050 438854
rect 271286 438618 271328 438854
rect 271008 438586 271328 438618
rect 301728 439174 302048 439206
rect 301728 438938 301770 439174
rect 302006 438938 302048 439174
rect 301728 438854 302048 438938
rect 301728 438618 301770 438854
rect 302006 438618 302048 438854
rect 301728 438586 302048 438618
rect 332448 439174 332768 439206
rect 332448 438938 332490 439174
rect 332726 438938 332768 439174
rect 332448 438854 332768 438938
rect 332448 438618 332490 438854
rect 332726 438618 332768 438854
rect 332448 438586 332768 438618
rect 363168 439174 363488 439206
rect 363168 438938 363210 439174
rect 363446 438938 363488 439174
rect 363168 438854 363488 438938
rect 363168 438618 363210 438854
rect 363446 438618 363488 438854
rect 363168 438586 363488 438618
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 255648 435454 255968 435486
rect 255648 435218 255690 435454
rect 255926 435218 255968 435454
rect 255648 435134 255968 435218
rect 255648 434898 255690 435134
rect 255926 434898 255968 435134
rect 255648 434866 255968 434898
rect 286368 435454 286688 435486
rect 286368 435218 286410 435454
rect 286646 435218 286688 435454
rect 286368 435134 286688 435218
rect 286368 434898 286410 435134
rect 286646 434898 286688 435134
rect 286368 434866 286688 434898
rect 317088 435454 317408 435486
rect 317088 435218 317130 435454
rect 317366 435218 317408 435454
rect 317088 435134 317408 435218
rect 317088 434898 317130 435134
rect 317366 434898 317408 435134
rect 317088 434866 317408 434898
rect 347808 435454 348128 435486
rect 347808 435218 347850 435454
rect 348086 435218 348128 435454
rect 347808 435134 348128 435218
rect 347808 434898 347850 435134
rect 348086 434898 348128 435134
rect 347808 434866 348128 434898
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 271008 403174 271328 403206
rect 271008 402938 271050 403174
rect 271286 402938 271328 403174
rect 271008 402854 271328 402938
rect 271008 402618 271050 402854
rect 271286 402618 271328 402854
rect 271008 402586 271328 402618
rect 301728 403174 302048 403206
rect 301728 402938 301770 403174
rect 302006 402938 302048 403174
rect 301728 402854 302048 402938
rect 301728 402618 301770 402854
rect 302006 402618 302048 402854
rect 301728 402586 302048 402618
rect 332448 403174 332768 403206
rect 332448 402938 332490 403174
rect 332726 402938 332768 403174
rect 332448 402854 332768 402938
rect 332448 402618 332490 402854
rect 332726 402618 332768 402854
rect 332448 402586 332768 402618
rect 363168 403174 363488 403206
rect 363168 402938 363210 403174
rect 363446 402938 363488 403174
rect 363168 402854 363488 402938
rect 363168 402618 363210 402854
rect 363446 402618 363488 402854
rect 363168 402586 363488 402618
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 255648 399454 255968 399486
rect 255648 399218 255690 399454
rect 255926 399218 255968 399454
rect 255648 399134 255968 399218
rect 255648 398898 255690 399134
rect 255926 398898 255968 399134
rect 255648 398866 255968 398898
rect 286368 399454 286688 399486
rect 286368 399218 286410 399454
rect 286646 399218 286688 399454
rect 286368 399134 286688 399218
rect 286368 398898 286410 399134
rect 286646 398898 286688 399134
rect 286368 398866 286688 398898
rect 317088 399454 317408 399486
rect 317088 399218 317130 399454
rect 317366 399218 317408 399454
rect 317088 399134 317408 399218
rect 317088 398898 317130 399134
rect 317366 398898 317408 399134
rect 317088 398866 317408 398898
rect 347808 399454 348128 399486
rect 347808 399218 347850 399454
rect 348086 399218 348128 399454
rect 347808 399134 348128 399218
rect 347808 398898 347850 399134
rect 348086 398898 348128 399134
rect 347808 398866 348128 398898
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 271008 367174 271328 367206
rect 271008 366938 271050 367174
rect 271286 366938 271328 367174
rect 271008 366854 271328 366938
rect 271008 366618 271050 366854
rect 271286 366618 271328 366854
rect 271008 366586 271328 366618
rect 301728 367174 302048 367206
rect 301728 366938 301770 367174
rect 302006 366938 302048 367174
rect 301728 366854 302048 366938
rect 301728 366618 301770 366854
rect 302006 366618 302048 366854
rect 301728 366586 302048 366618
rect 332448 367174 332768 367206
rect 332448 366938 332490 367174
rect 332726 366938 332768 367174
rect 332448 366854 332768 366938
rect 332448 366618 332490 366854
rect 332726 366618 332768 366854
rect 332448 366586 332768 366618
rect 363168 367174 363488 367206
rect 363168 366938 363210 367174
rect 363446 366938 363488 367174
rect 363168 366854 363488 366938
rect 363168 366618 363210 366854
rect 363446 366618 363488 366854
rect 363168 366586 363488 366618
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 255648 363454 255968 363486
rect 255648 363218 255690 363454
rect 255926 363218 255968 363454
rect 255648 363134 255968 363218
rect 255648 362898 255690 363134
rect 255926 362898 255968 363134
rect 255648 362866 255968 362898
rect 286368 363454 286688 363486
rect 286368 363218 286410 363454
rect 286646 363218 286688 363454
rect 286368 363134 286688 363218
rect 286368 362898 286410 363134
rect 286646 362898 286688 363134
rect 286368 362866 286688 362898
rect 317088 363454 317408 363486
rect 317088 363218 317130 363454
rect 317366 363218 317408 363454
rect 317088 363134 317408 363218
rect 317088 362898 317130 363134
rect 317366 362898 317408 363134
rect 317088 362866 317408 362898
rect 347808 363454 348128 363486
rect 347808 363218 347850 363454
rect 348086 363218 348128 363454
rect 347808 363134 348128 363218
rect 347808 362898 347850 363134
rect 348086 362898 348128 363134
rect 347808 362866 348128 362898
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 271008 331174 271328 331206
rect 271008 330938 271050 331174
rect 271286 330938 271328 331174
rect 271008 330854 271328 330938
rect 271008 330618 271050 330854
rect 271286 330618 271328 330854
rect 271008 330586 271328 330618
rect 301728 331174 302048 331206
rect 301728 330938 301770 331174
rect 302006 330938 302048 331174
rect 301728 330854 302048 330938
rect 301728 330618 301770 330854
rect 302006 330618 302048 330854
rect 301728 330586 302048 330618
rect 332448 331174 332768 331206
rect 332448 330938 332490 331174
rect 332726 330938 332768 331174
rect 332448 330854 332768 330938
rect 332448 330618 332490 330854
rect 332726 330618 332768 330854
rect 332448 330586 332768 330618
rect 363168 331174 363488 331206
rect 363168 330938 363210 331174
rect 363446 330938 363488 331174
rect 363168 330854 363488 330938
rect 363168 330618 363210 330854
rect 363446 330618 363488 330854
rect 363168 330586 363488 330618
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 255648 327454 255968 327486
rect 255648 327218 255690 327454
rect 255926 327218 255968 327454
rect 255648 327134 255968 327218
rect 255648 326898 255690 327134
rect 255926 326898 255968 327134
rect 255648 326866 255968 326898
rect 286368 327454 286688 327486
rect 286368 327218 286410 327454
rect 286646 327218 286688 327454
rect 286368 327134 286688 327218
rect 286368 326898 286410 327134
rect 286646 326898 286688 327134
rect 286368 326866 286688 326898
rect 317088 327454 317408 327486
rect 317088 327218 317130 327454
rect 317366 327218 317408 327454
rect 317088 327134 317408 327218
rect 317088 326898 317130 327134
rect 317366 326898 317408 327134
rect 317088 326866 317408 326898
rect 347808 327454 348128 327486
rect 347808 327218 347850 327454
rect 348086 327218 348128 327454
rect 347808 327134 348128 327218
rect 347808 326898 347850 327134
rect 348086 326898 348128 327134
rect 347808 326866 348128 326898
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 271008 295174 271328 295206
rect 271008 294938 271050 295174
rect 271286 294938 271328 295174
rect 271008 294854 271328 294938
rect 271008 294618 271050 294854
rect 271286 294618 271328 294854
rect 271008 294586 271328 294618
rect 301728 295174 302048 295206
rect 301728 294938 301770 295174
rect 302006 294938 302048 295174
rect 301728 294854 302048 294938
rect 301728 294618 301770 294854
rect 302006 294618 302048 294854
rect 301728 294586 302048 294618
rect 332448 295174 332768 295206
rect 332448 294938 332490 295174
rect 332726 294938 332768 295174
rect 332448 294854 332768 294938
rect 332448 294618 332490 294854
rect 332726 294618 332768 294854
rect 332448 294586 332768 294618
rect 363168 295174 363488 295206
rect 363168 294938 363210 295174
rect 363446 294938 363488 295174
rect 363168 294854 363488 294938
rect 363168 294618 363210 294854
rect 363446 294618 363488 294854
rect 363168 294586 363488 294618
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 255648 291454 255968 291486
rect 255648 291218 255690 291454
rect 255926 291218 255968 291454
rect 255648 291134 255968 291218
rect 255648 290898 255690 291134
rect 255926 290898 255968 291134
rect 255648 290866 255968 290898
rect 286368 291454 286688 291486
rect 286368 291218 286410 291454
rect 286646 291218 286688 291454
rect 286368 291134 286688 291218
rect 286368 290898 286410 291134
rect 286646 290898 286688 291134
rect 286368 290866 286688 290898
rect 317088 291454 317408 291486
rect 317088 291218 317130 291454
rect 317366 291218 317408 291454
rect 317088 291134 317408 291218
rect 317088 290898 317130 291134
rect 317366 290898 317408 291134
rect 317088 290866 317408 290898
rect 347808 291454 348128 291486
rect 347808 291218 347850 291454
rect 348086 291218 348128 291454
rect 347808 291134 348128 291218
rect 347808 290898 347850 291134
rect 348086 290898 348128 291134
rect 347808 290866 348128 290898
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 271008 259174 271328 259206
rect 271008 258938 271050 259174
rect 271286 258938 271328 259174
rect 271008 258854 271328 258938
rect 271008 258618 271050 258854
rect 271286 258618 271328 258854
rect 271008 258586 271328 258618
rect 301728 259174 302048 259206
rect 301728 258938 301770 259174
rect 302006 258938 302048 259174
rect 301728 258854 302048 258938
rect 301728 258618 301770 258854
rect 302006 258618 302048 258854
rect 301728 258586 302048 258618
rect 332448 259174 332768 259206
rect 332448 258938 332490 259174
rect 332726 258938 332768 259174
rect 332448 258854 332768 258938
rect 332448 258618 332490 258854
rect 332726 258618 332768 258854
rect 332448 258586 332768 258618
rect 363168 259174 363488 259206
rect 363168 258938 363210 259174
rect 363446 258938 363488 259174
rect 363168 258854 363488 258938
rect 363168 258618 363210 258854
rect 363446 258618 363488 258854
rect 363168 258586 363488 258618
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 255648 255454 255968 255486
rect 255648 255218 255690 255454
rect 255926 255218 255968 255454
rect 255648 255134 255968 255218
rect 255648 254898 255690 255134
rect 255926 254898 255968 255134
rect 255648 254866 255968 254898
rect 286368 255454 286688 255486
rect 286368 255218 286410 255454
rect 286646 255218 286688 255454
rect 286368 255134 286688 255218
rect 286368 254898 286410 255134
rect 286646 254898 286688 255134
rect 286368 254866 286688 254898
rect 317088 255454 317408 255486
rect 317088 255218 317130 255454
rect 317366 255218 317408 255454
rect 317088 255134 317408 255218
rect 317088 254898 317130 255134
rect 317366 254898 317408 255134
rect 317088 254866 317408 254898
rect 347808 255454 348128 255486
rect 347808 255218 347850 255454
rect 348086 255218 348128 255454
rect 347808 255134 348128 255218
rect 347808 254898 347850 255134
rect 348086 254898 348128 255134
rect 347808 254866 348128 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 223174 258134 249743
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 226894 261854 249743
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 230614 265574 249743
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 234334 269294 249743
rect 268674 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 269294 234334
rect 268674 234014 269294 234098
rect 268674 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 269294 234014
rect 268674 198334 269294 233778
rect 268674 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 269294 198334
rect 268674 198014 269294 198098
rect 268674 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 269294 198014
rect 268674 162334 269294 197778
rect 268674 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 269294 162334
rect 268674 162014 269294 162098
rect 268674 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 269294 162014
rect 268674 126334 269294 161778
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 268674 90334 269294 125778
rect 268674 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 269294 90334
rect 268674 90014 269294 90098
rect 268674 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 269294 90014
rect 268674 54334 269294 89778
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 238054 273014 249743
rect 272394 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 273014 238054
rect 272394 237734 273014 237818
rect 272394 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 273014 237734
rect 272394 202054 273014 237498
rect 272394 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 273014 202054
rect 272394 201734 273014 201818
rect 272394 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 273014 201734
rect 272394 166054 273014 201498
rect 272394 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 273014 166054
rect 272394 165734 273014 165818
rect 272394 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 273014 165734
rect 272394 130054 273014 165498
rect 272394 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 273014 130054
rect 272394 129734 273014 129818
rect 272394 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 273014 129734
rect 272394 94054 273014 129498
rect 272394 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 273014 94054
rect 272394 93734 273014 93818
rect 272394 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 273014 93734
rect 272394 58054 273014 93498
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 241774 276734 249743
rect 276114 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 276734 241774
rect 276114 241454 276734 241538
rect 276114 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 276734 241454
rect 276114 205774 276734 241218
rect 276114 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 276734 205774
rect 276114 205454 276734 205538
rect 276114 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 276734 205454
rect 276114 169774 276734 205218
rect 276114 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 276734 169774
rect 276114 169454 276734 169538
rect 276114 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 276734 169454
rect 276114 133774 276734 169218
rect 276114 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 276734 133774
rect 276114 133454 276734 133538
rect 276114 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 276734 133454
rect 276114 97774 276734 133218
rect 276114 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 276734 97774
rect 276114 97454 276734 97538
rect 276114 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 276734 97454
rect 276114 61774 276734 97218
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 276114 25774 276734 61218
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 245494 280454 249743
rect 279834 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 280454 245494
rect 279834 245174 280454 245258
rect 279834 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 280454 245174
rect 279834 209494 280454 244938
rect 279834 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 280454 209494
rect 279834 209174 280454 209258
rect 279834 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 280454 209174
rect 279834 173494 280454 208938
rect 279834 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 280454 173494
rect 279834 173174 280454 173258
rect 279834 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 280454 173174
rect 279834 137494 280454 172938
rect 279834 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 280454 137494
rect 279834 137174 280454 137258
rect 279834 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 280454 137174
rect 279834 101494 280454 136938
rect 279834 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 280454 101494
rect 279834 101174 280454 101258
rect 279834 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 280454 101174
rect 279834 65494 280454 100938
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 279834 29494 280454 64938
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 219454 290414 249743
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 223174 294134 249743
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 226894 297854 249743
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 230614 301574 249743
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 234334 305294 249743
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 304674 198334 305294 233778
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 304674 162334 305294 197778
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304674 90334 305294 125778
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 304674 54334 305294 89778
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 238054 309014 249743
rect 308394 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 309014 238054
rect 308394 237734 309014 237818
rect 308394 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 309014 237734
rect 308394 202054 309014 237498
rect 308394 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 309014 202054
rect 308394 201734 309014 201818
rect 308394 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 309014 201734
rect 308394 166054 309014 201498
rect 308394 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 309014 166054
rect 308394 165734 309014 165818
rect 308394 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 309014 165734
rect 308394 130054 309014 165498
rect 308394 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 309014 130054
rect 308394 129734 309014 129818
rect 308394 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 309014 129734
rect 308394 94054 309014 129498
rect 308394 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 309014 94054
rect 308394 93734 309014 93818
rect 308394 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 309014 93734
rect 308394 58054 309014 93498
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 241774 312734 249743
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 312114 205774 312734 241218
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 312114 169774 312734 205218
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 312114 133774 312734 169218
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 312114 97774 312734 133218
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 312114 61774 312734 97218
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 312114 25774 312734 61218
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 245494 316454 249743
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 101494 316454 136938
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 315834 65494 316454 100938
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 219454 326414 249743
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 223174 330134 249743
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 226894 333854 249743
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 230614 337574 249743
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 234334 341294 249743
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 340674 162334 341294 197778
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 340674 126334 341294 161778
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 90334 341294 125778
rect 340674 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 341294 90334
rect 340674 90014 341294 90098
rect 340674 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 341294 90014
rect 340674 54334 341294 89778
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 238054 345014 249743
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 344394 166054 345014 201498
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 344394 130054 345014 165498
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 344394 94054 345014 129498
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 344394 58054 345014 93498
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 241774 348734 249743
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 97774 348734 133218
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 245494 352454 249743
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351834 101494 352454 136938
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 219454 362414 249743
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 223174 366134 249743
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 378528 435454 378848 435486
rect 378528 435218 378570 435454
rect 378806 435218 378848 435454
rect 378528 435134 378848 435218
rect 378528 434898 378570 435134
rect 378806 434898 378848 435134
rect 378528 434866 378848 434898
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 378528 399454 378848 399486
rect 378528 399218 378570 399454
rect 378806 399218 378848 399454
rect 378528 399134 378848 399218
rect 378528 398898 378570 399134
rect 378806 398898 378848 399134
rect 378528 398866 378848 398898
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 378528 363454 378848 363486
rect 378528 363218 378570 363454
rect 378806 363218 378848 363454
rect 378528 363134 378848 363218
rect 378528 362898 378570 363134
rect 378806 362898 378848 363134
rect 378528 362866 378848 362898
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 378528 327454 378848 327486
rect 378528 327218 378570 327454
rect 378806 327218 378848 327454
rect 378528 327134 378848 327218
rect 378528 326898 378570 327134
rect 378806 326898 378848 327134
rect 378528 326866 378848 326898
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 378528 291454 378848 291486
rect 378528 291218 378570 291454
rect 378806 291218 378848 291454
rect 378528 291134 378848 291218
rect 378528 290898 378570 291134
rect 378806 290898 378848 291134
rect 378528 290866 378848 290898
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 378528 255454 378848 255486
rect 378528 255218 378570 255454
rect 378806 255218 378848 255454
rect 378528 255134 378848 255218
rect 378528 254898 378570 255134
rect 378806 254898 378848 255134
rect 378528 254866 378848 254898
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 389219 449716 389285 449717
rect 389219 449652 389220 449716
rect 389284 449652 389285 449716
rect 389219 449651 389285 449652
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 389222 48109 389282 449651
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 389219 48108 389285 48109
rect 389219 48044 389220 48108
rect 389284 48044 389285 48108
rect 389219 48043 389285 48044
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 585244 420734 601218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 585244 424454 604938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 585244 434414 614898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 585244 438134 618618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 585244 441854 586338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 585244 445574 590058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 585244 449294 593778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 585244 453014 597498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 585244 456734 601218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 641494 460454 676938
rect 459834 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 460454 641494
rect 459834 641174 460454 641258
rect 459834 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 460454 641174
rect 459834 605494 460454 640938
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 459834 585244 460454 604938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 585244 470414 614898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 585244 474134 618618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 585244 477854 586338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 585244 481574 590058
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484674 630334 485294 665778
rect 484674 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 485294 630334
rect 484674 630014 485294 630098
rect 484674 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 485294 630014
rect 484674 594334 485294 629778
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 585244 485294 593778
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 634054 489014 669498
rect 488394 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 489014 634054
rect 488394 633734 489014 633818
rect 488394 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 489014 633734
rect 488394 598054 489014 633498
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 585244 489014 597498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 637774 492734 673218
rect 492114 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 492734 637774
rect 492114 637454 492734 637538
rect 492114 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 492734 637454
rect 492114 601774 492734 637218
rect 492114 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 492734 601774
rect 492114 601454 492734 601538
rect 492114 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 492734 601454
rect 492114 585244 492734 601218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 641494 496454 676938
rect 495834 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 496454 641494
rect 495834 641174 496454 641258
rect 495834 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 496454 641174
rect 495834 605494 496454 640938
rect 495834 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 496454 605494
rect 495834 605174 496454 605258
rect 495834 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 496454 605174
rect 495834 585244 496454 604938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 585244 506414 614898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 585244 510134 618618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 585244 513854 586338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 585244 517574 590058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 585244 521294 593778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 585244 525014 597498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 585244 528734 601218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 585244 532454 604938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 585244 542414 614898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 585244 546134 618618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 585244 549854 586338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 585244 553574 590058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 585244 557294 593778
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 550955 585172 551021 585173
rect 550955 585108 550956 585172
rect 551020 585108 551021 585172
rect 550955 585107 551021 585108
rect 550958 583810 551018 585107
rect 550840 583750 551018 583810
rect 550840 583202 550900 583750
rect 420272 582929 420620 583036
rect 420272 582693 420328 582929
rect 420564 582693 420620 582929
rect 420272 582586 420620 582693
rect 556000 582929 556348 583036
rect 556000 582693 556056 582929
rect 556292 582693 556348 582929
rect 556000 582586 556348 582693
rect 420952 579454 421300 579486
rect 420952 579218 421008 579454
rect 421244 579218 421300 579454
rect 420952 579134 421300 579218
rect 420952 578898 421008 579134
rect 421244 578898 421300 579134
rect 420952 578866 421300 578898
rect 555320 579454 555668 579486
rect 555320 579218 555376 579454
rect 555612 579218 555668 579454
rect 555320 579134 555668 579218
rect 555320 578898 555376 579134
rect 555612 578898 555668 579134
rect 555320 578866 555668 578898
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 420272 547174 420620 547206
rect 420272 546938 420328 547174
rect 420564 546938 420620 547174
rect 420272 546854 420620 546938
rect 420272 546618 420328 546854
rect 420564 546618 420620 546854
rect 420272 546586 420620 546618
rect 556000 547174 556348 547206
rect 556000 546938 556056 547174
rect 556292 546938 556348 547174
rect 556000 546854 556348 546938
rect 556000 546618 556056 546854
rect 556292 546618 556348 546854
rect 556000 546586 556348 546618
rect 420952 543454 421300 543486
rect 420952 543218 421008 543454
rect 421244 543218 421300 543454
rect 420952 543134 421300 543218
rect 420952 542898 421008 543134
rect 421244 542898 421300 543134
rect 420952 542866 421300 542898
rect 555320 543454 555668 543486
rect 555320 543218 555376 543454
rect 555612 543218 555668 543454
rect 555320 543134 555668 543218
rect 555320 542898 555376 543134
rect 555612 542898 555668 543134
rect 555320 542866 555668 542898
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 420272 511174 420620 511206
rect 420272 510938 420328 511174
rect 420564 510938 420620 511174
rect 420272 510854 420620 510938
rect 420272 510618 420328 510854
rect 420564 510618 420620 510854
rect 420272 510586 420620 510618
rect 556000 511174 556348 511206
rect 556000 510938 556056 511174
rect 556292 510938 556348 511174
rect 556000 510854 556348 510938
rect 556000 510618 556056 510854
rect 556292 510618 556348 510854
rect 556000 510586 556348 510618
rect 420952 507454 421300 507486
rect 420952 507218 421008 507454
rect 421244 507218 421300 507454
rect 420952 507134 421300 507218
rect 420952 506898 421008 507134
rect 421244 506898 421300 507134
rect 420952 506866 421300 506898
rect 555320 507454 555668 507486
rect 555320 507218 555376 507454
rect 555612 507218 555668 507454
rect 555320 507134 555668 507218
rect 555320 506898 555376 507134
rect 555612 506898 555668 507134
rect 555320 506866 555668 506898
rect 436056 499590 436116 500106
rect 437144 499590 437204 500106
rect 436056 499530 436202 499590
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 420114 493774 420734 498064
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 418659 462772 418725 462773
rect 418659 462708 418660 462772
rect 418724 462708 418725 462772
rect 418659 462707 418725 462708
rect 418107 454612 418173 454613
rect 418107 454548 418108 454612
rect 418172 454548 418173 454612
rect 418107 454547 418173 454548
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 415899 450260 415965 450261
rect 415899 450196 415900 450260
rect 415964 450196 415965 450260
rect 415899 450195 415965 450196
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 306334 413294 341778
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 415902 47701 415962 450195
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 417923 359956 417989 359957
rect 417923 359892 417924 359956
rect 417988 359892 417989 359956
rect 417923 359891 417989 359892
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 416394 310054 417014 345498
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 417739 278764 417805 278765
rect 417739 278700 417740 278764
rect 417804 278700 417805 278764
rect 417739 278699 417805 278700
rect 417742 278221 417802 278699
rect 417739 278220 417805 278221
rect 417739 278156 417740 278220
rect 417804 278156 417805 278220
rect 417739 278155 417805 278156
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 417555 260812 417621 260813
rect 417555 260748 417556 260812
rect 417620 260748 417621 260812
rect 417555 260747 417621 260748
rect 417558 259997 417618 260747
rect 417555 259996 417621 259997
rect 417555 259932 417556 259996
rect 417620 259932 417621 259996
rect 417555 259931 417621 259932
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 130054 417014 165498
rect 417558 160037 417618 259931
rect 417742 178261 417802 278155
rect 417926 260813 417986 359891
rect 417923 260812 417989 260813
rect 417923 260748 417924 260812
rect 417988 260748 417989 260812
rect 417923 260747 417989 260748
rect 418110 249525 418170 454547
rect 418107 249524 418173 249525
rect 418107 249460 418108 249524
rect 418172 249460 418173 249524
rect 418107 249459 418173 249460
rect 417923 179484 417989 179485
rect 417923 179420 417924 179484
rect 417988 179420 417989 179484
rect 417923 179419 417989 179420
rect 417739 178260 417805 178261
rect 417739 178196 417740 178260
rect 417804 178196 417805 178260
rect 417739 178195 417805 178196
rect 417555 160036 417621 160037
rect 417555 159972 417556 160036
rect 417620 159972 417621 160036
rect 417555 159971 417621 159972
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 417558 59941 417618 159971
rect 417742 78165 417802 178195
rect 417926 79933 417986 179419
rect 417923 79932 417989 79933
rect 417923 79868 417924 79932
rect 417988 79868 417989 79932
rect 417923 79867 417989 79868
rect 417739 78164 417805 78165
rect 417739 78100 417740 78164
rect 417804 78100 417805 78164
rect 417739 78099 417805 78100
rect 417555 59940 417621 59941
rect 417555 59876 417556 59940
rect 417620 59876 417621 59940
rect 417555 59875 417621 59876
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 415899 47700 415965 47701
rect 415899 47636 415900 47700
rect 415964 47636 415965 47700
rect 415899 47635 415965 47636
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 57498
rect 418662 49197 418722 462707
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 418843 450532 418909 450533
rect 418843 450468 418844 450532
rect 418908 450468 418909 450532
rect 418843 450467 418909 450468
rect 418846 249525 418906 450467
rect 420114 435244 420734 457218
rect 423834 497494 424454 498064
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 435244 424454 460938
rect 433794 471454 434414 498064
rect 436142 497181 436202 499530
rect 437062 499530 437204 499590
rect 438232 499590 438292 500106
rect 439592 499590 439652 500106
rect 440544 499590 440604 500106
rect 441768 499590 441828 500106
rect 438232 499530 438410 499590
rect 439592 499530 439698 499590
rect 440544 499530 440618 499590
rect 437062 497317 437122 499530
rect 437059 497316 437125 497317
rect 437059 497252 437060 497316
rect 437124 497252 437125 497316
rect 437059 497251 437125 497252
rect 436139 497180 436205 497181
rect 436139 497116 436140 497180
rect 436204 497116 436205 497180
rect 436139 497115 436205 497116
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435244 434414 470898
rect 437514 475174 438134 498064
rect 438350 496909 438410 499530
rect 439638 496909 439698 499530
rect 440558 496909 440618 499530
rect 441662 499530 441828 499590
rect 443128 499590 443188 500106
rect 444216 499590 444276 500106
rect 445440 499590 445500 500106
rect 446528 499590 446588 500106
rect 447616 499590 447676 500106
rect 448296 499590 448356 500106
rect 448704 499590 448764 500106
rect 450064 499590 450124 500106
rect 450744 499590 450804 500106
rect 443128 499530 443194 499590
rect 444216 499530 444298 499590
rect 441662 498133 441722 499530
rect 441659 498132 441725 498133
rect 441659 498068 441660 498132
rect 441724 498068 441725 498132
rect 441659 498067 441725 498068
rect 438347 496908 438413 496909
rect 438347 496844 438348 496908
rect 438412 496844 438413 496908
rect 438347 496843 438413 496844
rect 439635 496908 439701 496909
rect 439635 496844 439636 496908
rect 439700 496844 439701 496908
rect 439635 496843 439701 496844
rect 440555 496908 440621 496909
rect 440555 496844 440556 496908
rect 440620 496844 440621 496908
rect 440555 496843 440621 496844
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 435244 438134 438618
rect 441234 478894 441854 497940
rect 443134 496909 443194 499530
rect 444238 497045 444298 499530
rect 445342 499530 445500 499590
rect 446446 499530 446588 499590
rect 447550 499530 447676 499590
rect 448286 499530 448356 499590
rect 448654 499530 448764 499590
rect 449942 499530 450124 499590
rect 450678 499530 450804 499590
rect 445342 498133 445402 499530
rect 445339 498132 445405 498133
rect 445339 498068 445340 498132
rect 445404 498068 445405 498132
rect 445339 498067 445405 498068
rect 444235 497044 444301 497045
rect 444235 496980 444236 497044
rect 444300 496980 444301 497044
rect 444235 496979 444301 496980
rect 443131 496908 443197 496909
rect 443131 496844 443132 496908
rect 443196 496844 443197 496908
rect 443131 496843 443197 496844
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 435244 441854 442338
rect 444954 482614 445574 497940
rect 446446 496909 446506 499530
rect 447550 496909 447610 499530
rect 448286 497045 448346 499530
rect 448654 498133 448714 499530
rect 448651 498132 448717 498133
rect 448651 498068 448652 498132
rect 448716 498068 448717 498132
rect 448651 498067 448717 498068
rect 448283 497044 448349 497045
rect 448283 496980 448284 497044
rect 448348 496980 448349 497044
rect 448283 496979 448349 496980
rect 446443 496908 446509 496909
rect 446443 496844 446444 496908
rect 446508 496844 446509 496908
rect 446443 496843 446509 496844
rect 447547 496908 447613 496909
rect 447547 496844 447548 496908
rect 447612 496844 447613 496908
rect 447547 496843 447613 496844
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 435244 445574 446058
rect 448674 486334 449294 497940
rect 449942 496909 450002 499530
rect 450678 497045 450738 499530
rect 451288 499490 451348 500106
rect 452376 499590 452436 500106
rect 453464 499590 453524 500106
rect 451046 499430 451348 499490
rect 452334 499530 452436 499590
rect 453438 499530 453524 499590
rect 453600 499590 453660 500106
rect 454552 499590 454612 500106
rect 453600 499530 453682 499590
rect 450675 497044 450741 497045
rect 450675 496980 450676 497044
rect 450740 496980 450741 497044
rect 450675 496979 450741 496980
rect 451046 496909 451106 499430
rect 452334 498133 452394 499530
rect 452331 498132 452397 498133
rect 452331 498068 452332 498132
rect 452396 498068 452397 498132
rect 452331 498067 452397 498068
rect 449939 496908 450005 496909
rect 449939 496844 449940 496908
rect 450004 496844 450005 496908
rect 449939 496843 450005 496844
rect 451043 496908 451109 496909
rect 451043 496844 451044 496908
rect 451108 496844 451109 496908
rect 451043 496843 451109 496844
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 435244 449294 449778
rect 452394 490054 453014 497940
rect 453438 497589 453498 499530
rect 453435 497588 453501 497589
rect 453435 497524 453436 497588
rect 453500 497524 453501 497588
rect 453435 497523 453501 497524
rect 453622 496909 453682 499530
rect 454542 499530 454612 499590
rect 454542 496909 454602 499530
rect 455912 499490 455972 500106
rect 456048 499590 456108 500106
rect 457000 499590 457060 500106
rect 458088 499590 458148 500106
rect 458496 499590 458556 500106
rect 459448 499590 459508 500106
rect 460672 499590 460732 500106
rect 461080 499590 461140 500106
rect 456048 499530 456258 499590
rect 455830 499430 455972 499490
rect 455830 497181 455890 499430
rect 456198 498133 456258 499530
rect 456934 499530 457060 499590
rect 458038 499530 458148 499590
rect 458406 499530 458556 499590
rect 459326 499530 459508 499590
rect 460614 499530 460732 499590
rect 460982 499530 461140 499590
rect 463528 499590 463588 500106
rect 465976 499590 466036 500106
rect 463528 499530 463618 499590
rect 456195 498132 456261 498133
rect 456195 498068 456196 498132
rect 456260 498068 456261 498132
rect 456195 498067 456261 498068
rect 455827 497180 455893 497181
rect 455827 497116 455828 497180
rect 455892 497116 455893 497180
rect 455827 497115 455893 497116
rect 453619 496908 453685 496909
rect 453619 496844 453620 496908
rect 453684 496844 453685 496908
rect 453619 496843 453685 496844
rect 454539 496908 454605 496909
rect 454539 496844 454540 496908
rect 454604 496844 454605 496908
rect 454539 496843 454605 496844
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 435244 453014 453498
rect 456114 493774 456734 497940
rect 456934 497045 456994 499530
rect 456931 497044 456997 497045
rect 456931 496980 456932 497044
rect 456996 496980 456997 497044
rect 456931 496979 456997 496980
rect 458038 496909 458098 499530
rect 458406 496909 458466 499530
rect 459326 497045 459386 499530
rect 459834 497494 460454 498064
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459323 497044 459389 497045
rect 459323 496980 459324 497044
rect 459388 496980 459389 497044
rect 459323 496979 459389 496980
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 460614 497045 460674 499530
rect 460611 497044 460677 497045
rect 460611 496980 460612 497044
rect 460676 496980 460677 497044
rect 460611 496979 460677 496980
rect 458035 496908 458101 496909
rect 458035 496844 458036 496908
rect 458100 496844 458101 496908
rect 458035 496843 458101 496844
rect 458403 496908 458469 496909
rect 458403 496844 458404 496908
rect 458468 496844 458469 496908
rect 458403 496843 458469 496844
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 435244 456734 457218
rect 459834 461494 460454 496938
rect 460982 496909 461042 499530
rect 463558 496909 463618 499530
rect 465950 499530 466036 499590
rect 468288 499590 468348 500106
rect 471008 499590 471068 500106
rect 473592 499590 473652 500106
rect 468288 499530 468402 499590
rect 465950 496909 466010 499530
rect 468342 496909 468402 499530
rect 470918 499530 471068 499590
rect 473494 499530 473652 499590
rect 476040 499590 476100 500106
rect 478488 499590 478548 500106
rect 480936 499590 480996 500106
rect 483520 499590 483580 500106
rect 476040 499530 476130 499590
rect 460979 496908 461045 496909
rect 460979 496844 460980 496908
rect 461044 496844 461045 496908
rect 460979 496843 461045 496844
rect 463555 496908 463621 496909
rect 463555 496844 463556 496908
rect 463620 496844 463621 496908
rect 463555 496843 463621 496844
rect 465947 496908 466013 496909
rect 465947 496844 465948 496908
rect 466012 496844 466013 496908
rect 465947 496843 466013 496844
rect 468339 496908 468405 496909
rect 468339 496844 468340 496908
rect 468404 496844 468405 496908
rect 468339 496843 468405 496844
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 435244 460454 460938
rect 469794 471454 470414 497940
rect 470918 497045 470978 499530
rect 473494 498133 473554 499530
rect 473491 498132 473557 498133
rect 473491 498068 473492 498132
rect 473556 498068 473557 498132
rect 473491 498067 473557 498068
rect 470915 497044 470981 497045
rect 470915 496980 470916 497044
rect 470980 496980 470981 497044
rect 470915 496979 470981 496980
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435244 470414 470898
rect 473514 475174 474134 497940
rect 476070 497045 476130 499530
rect 478462 499530 478548 499590
rect 480854 499530 480996 499590
rect 483430 499530 483580 499590
rect 485968 499590 486028 500106
rect 485968 499530 486066 499590
rect 476067 497044 476133 497045
rect 476067 496980 476068 497044
rect 476132 496980 476133 497044
rect 476067 496979 476133 496980
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 435244 474134 438618
rect 477234 478894 477854 498064
rect 478462 496909 478522 499530
rect 480854 498133 480914 499530
rect 480851 498132 480917 498133
rect 480851 498068 480852 498132
rect 480916 498068 480917 498132
rect 480851 498067 480917 498068
rect 478459 496908 478525 496909
rect 478459 496844 478460 496908
rect 478524 496844 478525 496908
rect 478459 496843 478525 496844
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 435244 477854 442338
rect 480954 482614 481574 497940
rect 483430 497181 483490 499530
rect 483427 497180 483493 497181
rect 483427 497116 483428 497180
rect 483492 497116 483493 497180
rect 483427 497115 483493 497116
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 435244 481574 446058
rect 484674 486334 485294 498064
rect 486006 497997 486066 499530
rect 486003 497996 486069 497997
rect 486003 497932 486004 497996
rect 486068 497932 486069 497996
rect 486003 497931 486069 497932
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 484674 435244 485294 449778
rect 488394 490054 489014 497940
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454054 489014 489498
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 488394 435244 489014 453498
rect 492114 493774 492734 498064
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 492114 435244 492734 457218
rect 495834 497494 496454 497940
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 435244 496454 460938
rect 505794 471454 506414 497940
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435244 506414 470898
rect 509514 475174 510134 498064
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 435244 510134 438618
rect 513234 478894 513854 497940
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 435244 513854 442338
rect 516954 482614 517574 498064
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 435244 517574 446058
rect 520674 486334 521294 497940
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 435244 521294 449778
rect 524394 490054 525014 498064
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 435244 525014 453498
rect 528114 493774 528734 498064
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 435244 528734 457218
rect 531834 497494 532454 498064
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 435244 532454 460938
rect 541794 471454 542414 498064
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435244 542414 470898
rect 545514 475174 546134 498064
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 435244 546134 438618
rect 549234 478894 549854 498064
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 435244 549854 442338
rect 552954 482614 553574 498064
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 435244 553574 446058
rect 556674 486334 557294 498064
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 435244 557294 449778
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 550837 433532 550903 433533
rect 550837 433468 550838 433532
rect 550902 433468 550903 433532
rect 550837 433467 550903 433468
rect 550840 433202 550900 433467
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 420272 403174 420620 403206
rect 420272 402938 420328 403174
rect 420564 402938 420620 403174
rect 420272 402854 420620 402938
rect 420272 402618 420328 402854
rect 420564 402618 420620 402854
rect 420272 402586 420620 402618
rect 556000 403174 556348 403206
rect 556000 402938 556056 403174
rect 556292 402938 556348 403174
rect 556000 402854 556348 402938
rect 556000 402618 556056 402854
rect 556292 402618 556348 402854
rect 556000 402586 556348 402618
rect 420952 399454 421300 399486
rect 420952 399218 421008 399454
rect 421244 399218 421300 399454
rect 420952 399134 421300 399218
rect 420952 398898 421008 399134
rect 421244 398898 421300 399134
rect 420952 398866 421300 398898
rect 555320 399454 555668 399486
rect 555320 399218 555376 399454
rect 555612 399218 555668 399454
rect 555320 399134 555668 399218
rect 555320 398898 555376 399134
rect 555612 398898 555668 399134
rect 555320 398866 555668 398898
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 420272 367174 420620 367206
rect 420272 366938 420328 367174
rect 420564 366938 420620 367174
rect 420272 366854 420620 366938
rect 420272 366618 420328 366854
rect 420564 366618 420620 366854
rect 420272 366586 420620 366618
rect 556000 367174 556348 367206
rect 556000 366938 556056 367174
rect 556292 366938 556348 367174
rect 556000 366854 556348 366938
rect 556000 366618 556056 366854
rect 556292 366618 556348 366854
rect 556000 366586 556348 366618
rect 420952 363454 421300 363486
rect 420952 363218 421008 363454
rect 421244 363218 421300 363454
rect 420952 363134 421300 363218
rect 420952 362898 421008 363134
rect 421244 362898 421300 363134
rect 420952 362866 421300 362898
rect 555320 363454 555668 363486
rect 555320 363218 555376 363454
rect 555612 363218 555668 363454
rect 555320 363134 555668 363218
rect 555320 362898 555376 363134
rect 555612 362898 555668 363134
rect 555320 362866 555668 362898
rect 436056 349890 436116 350106
rect 437144 349890 437204 350106
rect 438232 349890 438292 350106
rect 436056 349830 436202 349890
rect 419763 347852 419829 347853
rect 419763 347788 419764 347852
rect 419828 347788 419829 347852
rect 419763 347787 419829 347788
rect 419579 346900 419645 346901
rect 419579 346836 419580 346900
rect 419644 346836 419645 346900
rect 419579 346835 419645 346836
rect 418843 249524 418909 249525
rect 418843 249460 418844 249524
rect 418908 249460 418909 249524
rect 418843 249459 418909 249460
rect 419211 235924 419277 235925
rect 419211 235860 419212 235924
rect 419276 235860 419277 235924
rect 419211 235859 419277 235860
rect 419214 146845 419274 235859
rect 419582 235789 419642 346835
rect 419766 248430 419826 347787
rect 436142 347717 436202 349830
rect 437062 349830 437204 349890
rect 438166 349830 438292 349890
rect 439592 349890 439652 350106
rect 440544 349890 440604 350106
rect 441768 349890 441828 350106
rect 439592 349830 439698 349890
rect 440544 349830 440618 349890
rect 437062 347717 437122 349830
rect 438166 347717 438226 349830
rect 439638 347717 439698 349830
rect 440558 347717 440618 349830
rect 441662 349830 441828 349890
rect 443128 349890 443188 350106
rect 444216 349890 444276 350106
rect 445440 349890 445500 350106
rect 446528 349890 446588 350106
rect 447616 349890 447676 350106
rect 448296 349890 448356 350106
rect 448704 349890 448764 350106
rect 443128 349830 443194 349890
rect 444216 349830 444298 349890
rect 441662 347717 441722 349830
rect 443134 347717 443194 349830
rect 444238 347717 444298 349830
rect 445342 349830 445500 349890
rect 446446 349830 446588 349890
rect 447550 349830 447676 349890
rect 448286 349830 448356 349890
rect 448654 349830 448764 349890
rect 450064 349890 450124 350106
rect 450744 349890 450804 350106
rect 450064 349830 450186 349890
rect 445342 347717 445402 349830
rect 446446 347717 446506 349830
rect 447550 347717 447610 349830
rect 448286 347717 448346 349830
rect 448654 347717 448714 349830
rect 450126 347717 450186 349830
rect 450678 349830 450804 349890
rect 451288 349890 451348 350106
rect 451288 349830 451474 349890
rect 450678 347717 450738 349830
rect 451414 347717 451474 349830
rect 452376 349757 452436 350106
rect 453464 349890 453524 350106
rect 453438 349830 453524 349890
rect 453600 349890 453660 350106
rect 454552 349890 454612 350106
rect 455912 349890 455972 350106
rect 453600 349830 453682 349890
rect 452373 349756 452439 349757
rect 452373 349692 452374 349756
rect 452438 349692 452439 349756
rect 452373 349691 452439 349692
rect 453438 347717 453498 349830
rect 453622 347717 453682 349830
rect 454542 349830 454612 349890
rect 455830 349830 455972 349890
rect 456048 349890 456108 350106
rect 457000 349890 457060 350106
rect 458088 349890 458148 350106
rect 458496 349890 458556 350106
rect 456048 349830 456258 349890
rect 454542 347717 454602 349830
rect 455830 347717 455890 349830
rect 456198 347717 456258 349830
rect 456934 349830 457060 349890
rect 458038 349830 458148 349890
rect 458406 349830 458556 349890
rect 459448 349890 459508 350106
rect 460672 349890 460732 350106
rect 461080 349890 461140 350106
rect 459448 349830 459570 349890
rect 456934 347717 456994 349830
rect 458038 347717 458098 349830
rect 458406 347717 458466 349830
rect 459510 347717 459570 349830
rect 460614 349830 460732 349890
rect 460982 349830 461140 349890
rect 436139 347716 436205 347717
rect 436139 347652 436140 347716
rect 436204 347652 436205 347716
rect 436139 347651 436205 347652
rect 437059 347716 437125 347717
rect 437059 347652 437060 347716
rect 437124 347652 437125 347716
rect 437059 347651 437125 347652
rect 438163 347716 438229 347717
rect 438163 347652 438164 347716
rect 438228 347652 438229 347716
rect 438163 347651 438229 347652
rect 439635 347716 439701 347717
rect 439635 347652 439636 347716
rect 439700 347652 439701 347716
rect 439635 347651 439701 347652
rect 440555 347716 440621 347717
rect 440555 347652 440556 347716
rect 440620 347652 440621 347716
rect 440555 347651 440621 347652
rect 441659 347716 441725 347717
rect 441659 347652 441660 347716
rect 441724 347652 441725 347716
rect 441659 347651 441725 347652
rect 443131 347716 443197 347717
rect 443131 347652 443132 347716
rect 443196 347652 443197 347716
rect 443131 347651 443197 347652
rect 444235 347716 444301 347717
rect 444235 347652 444236 347716
rect 444300 347652 444301 347716
rect 444235 347651 444301 347652
rect 445339 347716 445405 347717
rect 445339 347652 445340 347716
rect 445404 347652 445405 347716
rect 445339 347651 445405 347652
rect 446443 347716 446509 347717
rect 446443 347652 446444 347716
rect 446508 347652 446509 347716
rect 446443 347651 446509 347652
rect 447547 347716 447613 347717
rect 447547 347652 447548 347716
rect 447612 347652 447613 347716
rect 447547 347651 447613 347652
rect 448283 347716 448349 347717
rect 448283 347652 448284 347716
rect 448348 347652 448349 347716
rect 448283 347651 448349 347652
rect 448651 347716 448717 347717
rect 448651 347652 448652 347716
rect 448716 347652 448717 347716
rect 448651 347651 448717 347652
rect 450123 347716 450189 347717
rect 450123 347652 450124 347716
rect 450188 347652 450189 347716
rect 450123 347651 450189 347652
rect 450675 347716 450741 347717
rect 450675 347652 450676 347716
rect 450740 347652 450741 347716
rect 450675 347651 450741 347652
rect 451411 347716 451477 347717
rect 451411 347652 451412 347716
rect 451476 347652 451477 347716
rect 451411 347651 451477 347652
rect 453435 347716 453501 347717
rect 453435 347652 453436 347716
rect 453500 347652 453501 347716
rect 453435 347651 453501 347652
rect 453619 347716 453685 347717
rect 453619 347652 453620 347716
rect 453684 347652 453685 347716
rect 453619 347651 453685 347652
rect 454539 347716 454605 347717
rect 454539 347652 454540 347716
rect 454604 347652 454605 347716
rect 454539 347651 454605 347652
rect 455827 347716 455893 347717
rect 455827 347652 455828 347716
rect 455892 347652 455893 347716
rect 455827 347651 455893 347652
rect 456195 347716 456261 347717
rect 456195 347652 456196 347716
rect 456260 347652 456261 347716
rect 456195 347651 456261 347652
rect 456931 347716 456997 347717
rect 456931 347652 456932 347716
rect 456996 347652 456997 347716
rect 456931 347651 456997 347652
rect 458035 347716 458101 347717
rect 458035 347652 458036 347716
rect 458100 347652 458101 347716
rect 458035 347651 458101 347652
rect 458403 347716 458469 347717
rect 458403 347652 458404 347716
rect 458468 347652 458469 347716
rect 458403 347651 458469 347652
rect 459507 347716 459573 347717
rect 459507 347652 459508 347716
rect 459572 347652 459573 347716
rect 459507 347651 459573 347652
rect 460614 347037 460674 349830
rect 460982 347717 461042 349830
rect 461760 349618 461820 350106
rect 462848 349618 462908 350106
rect 461718 349558 461820 349618
rect 462822 349558 462908 349618
rect 463528 349618 463588 350106
rect 463936 349618 463996 350106
rect 465296 349890 465356 350106
rect 463528 349558 463618 349618
rect 461718 347717 461778 349558
rect 462822 347717 462882 349558
rect 463558 347717 463618 349558
rect 463926 349558 463996 349618
rect 465214 349830 465356 349890
rect 463926 347717 463986 349558
rect 465214 347717 465274 349830
rect 465976 349618 466036 350106
rect 466384 349890 466444 350106
rect 465950 349558 466036 349618
rect 466318 349830 466444 349890
rect 460979 347716 461045 347717
rect 460979 347652 460980 347716
rect 461044 347652 461045 347716
rect 460979 347651 461045 347652
rect 461715 347716 461781 347717
rect 461715 347652 461716 347716
rect 461780 347652 461781 347716
rect 461715 347651 461781 347652
rect 462819 347716 462885 347717
rect 462819 347652 462820 347716
rect 462884 347652 462885 347716
rect 462819 347651 462885 347652
rect 463555 347716 463621 347717
rect 463555 347652 463556 347716
rect 463620 347652 463621 347716
rect 463555 347651 463621 347652
rect 463923 347716 463989 347717
rect 463923 347652 463924 347716
rect 463988 347652 463989 347716
rect 463923 347651 463989 347652
rect 465211 347716 465277 347717
rect 465211 347652 465212 347716
rect 465276 347652 465277 347716
rect 465211 347651 465277 347652
rect 465950 347037 466010 349558
rect 466318 347717 466378 349830
rect 467608 349618 467668 350106
rect 467606 349558 467668 349618
rect 468288 349618 468348 350106
rect 468696 349618 468756 350106
rect 469784 349618 469844 350106
rect 471008 349890 471068 350106
rect 470366 349830 471068 349890
rect 471144 349890 471204 350106
rect 472232 349890 472292 350106
rect 473320 349890 473380 350106
rect 473592 349890 473652 350106
rect 471144 349830 471346 349890
rect 468288 349558 468402 349618
rect 468696 349558 468770 349618
rect 469784 349558 469874 349618
rect 467606 347717 467666 349558
rect 466315 347716 466381 347717
rect 466315 347652 466316 347716
rect 466380 347652 466381 347716
rect 466315 347651 466381 347652
rect 467603 347716 467669 347717
rect 467603 347652 467604 347716
rect 467668 347652 467669 347716
rect 467603 347651 467669 347652
rect 468342 347581 468402 349558
rect 468710 347717 468770 349558
rect 469814 347717 469874 349558
rect 468707 347716 468773 347717
rect 468707 347652 468708 347716
rect 468772 347652 468773 347716
rect 468707 347651 468773 347652
rect 469811 347716 469877 347717
rect 469811 347652 469812 347716
rect 469876 347652 469877 347716
rect 469811 347651 469877 347652
rect 470366 347581 470426 349830
rect 471286 347717 471346 349830
rect 472206 349830 472292 349890
rect 473310 349830 473380 349890
rect 473494 349830 473652 349890
rect 474408 349890 474468 350106
rect 475768 349890 475828 350106
rect 474408 349830 474474 349890
rect 472206 347717 472266 349830
rect 473310 347717 473370 349830
rect 471283 347716 471349 347717
rect 471283 347652 471284 347716
rect 471348 347652 471349 347716
rect 471283 347651 471349 347652
rect 472203 347716 472269 347717
rect 472203 347652 472204 347716
rect 472268 347652 472269 347716
rect 472203 347651 472269 347652
rect 473307 347716 473373 347717
rect 473307 347652 473308 347716
rect 473372 347652 473373 347716
rect 473307 347651 473373 347652
rect 468339 347580 468405 347581
rect 468339 347516 468340 347580
rect 468404 347516 468405 347580
rect 468339 347515 468405 347516
rect 470363 347580 470429 347581
rect 470363 347516 470364 347580
rect 470428 347516 470429 347580
rect 470363 347515 470429 347516
rect 473494 347445 473554 349830
rect 474414 347717 474474 349830
rect 475702 349830 475828 349890
rect 476040 349890 476100 350106
rect 476992 349890 477052 350106
rect 476040 349830 476130 349890
rect 475702 347717 475762 349830
rect 474411 347716 474477 347717
rect 474411 347652 474412 347716
rect 474476 347652 474477 347716
rect 474411 347651 474477 347652
rect 475699 347716 475765 347717
rect 475699 347652 475700 347716
rect 475764 347652 475765 347716
rect 475699 347651 475765 347652
rect 473491 347444 473557 347445
rect 473491 347380 473492 347444
rect 473556 347380 473557 347444
rect 473491 347379 473557 347380
rect 476070 347309 476130 349830
rect 476990 349830 477052 349890
rect 478080 349890 478140 350106
rect 478488 349893 478548 350106
rect 478485 349892 478551 349893
rect 478080 349830 478154 349890
rect 476990 347717 477050 349830
rect 478094 347717 478154 349830
rect 478485 349828 478486 349892
rect 478550 349828 478551 349892
rect 479168 349890 479228 350106
rect 480936 349890 480996 350106
rect 483520 349893 483580 350106
rect 485968 349893 486028 350106
rect 479168 349830 479258 349890
rect 478485 349827 478551 349828
rect 479198 347717 479258 349830
rect 480854 349830 480996 349890
rect 483517 349892 483583 349893
rect 480854 349213 480914 349830
rect 483517 349828 483518 349892
rect 483582 349828 483583 349892
rect 483517 349827 483583 349828
rect 485965 349892 486031 349893
rect 485965 349828 485966 349892
rect 486030 349828 486031 349892
rect 485965 349827 486031 349828
rect 488280 349757 488340 350106
rect 491000 349757 491060 350106
rect 493448 349890 493508 350106
rect 495896 349893 495956 350106
rect 493366 349830 493508 349890
rect 495893 349892 495959 349893
rect 488277 349756 488343 349757
rect 488277 349692 488278 349756
rect 488342 349692 488343 349756
rect 488277 349691 488343 349692
rect 490997 349756 491063 349757
rect 490997 349692 490998 349756
rect 491062 349692 491063 349756
rect 490997 349691 491063 349692
rect 480851 349212 480917 349213
rect 480851 349148 480852 349212
rect 480916 349148 480917 349212
rect 480851 349147 480917 349148
rect 476987 347716 477053 347717
rect 476987 347652 476988 347716
rect 477052 347652 477053 347716
rect 476987 347651 477053 347652
rect 478091 347716 478157 347717
rect 478091 347652 478092 347716
rect 478156 347652 478157 347716
rect 478091 347651 478157 347652
rect 479195 347716 479261 347717
rect 479195 347652 479196 347716
rect 479260 347652 479261 347716
rect 479195 347651 479261 347652
rect 476067 347308 476133 347309
rect 476067 347244 476068 347308
rect 476132 347244 476133 347308
rect 476067 347243 476133 347244
rect 493366 347173 493426 349830
rect 495893 349828 495894 349892
rect 495958 349828 495959 349892
rect 498480 349890 498540 350106
rect 500928 349890 500988 350106
rect 503512 349890 503572 350106
rect 498480 349830 498578 349890
rect 495893 349827 495959 349828
rect 498518 349077 498578 349830
rect 500910 349830 500988 349890
rect 503486 349830 503572 349890
rect 500910 349077 500970 349830
rect 503486 349077 503546 349830
rect 505960 349621 506020 350106
rect 508544 349757 508604 350106
rect 510992 349890 511052 350106
rect 513440 349890 513500 350106
rect 510992 349830 511090 349890
rect 508541 349756 508607 349757
rect 508541 349692 508542 349756
rect 508606 349692 508607 349756
rect 508541 349691 508607 349692
rect 505957 349620 506023 349621
rect 505957 349556 505958 349620
rect 506022 349556 506023 349620
rect 505957 349555 506023 349556
rect 511030 349077 511090 349830
rect 513422 349830 513500 349890
rect 498515 349076 498581 349077
rect 498515 349012 498516 349076
rect 498580 349012 498581 349076
rect 498515 349011 498581 349012
rect 500907 349076 500973 349077
rect 500907 349012 500908 349076
rect 500972 349012 500973 349076
rect 500907 349011 500973 349012
rect 503483 349076 503549 349077
rect 503483 349012 503484 349076
rect 503548 349012 503549 349076
rect 503483 349011 503549 349012
rect 511027 349076 511093 349077
rect 511027 349012 511028 349076
rect 511092 349012 511093 349076
rect 511027 349011 511093 349012
rect 513422 347717 513482 349830
rect 515888 349621 515948 350106
rect 518472 349890 518532 350106
rect 518390 349830 518532 349890
rect 515885 349620 515951 349621
rect 515885 349556 515886 349620
rect 515950 349556 515951 349620
rect 515885 349555 515951 349556
rect 518390 347717 518450 349830
rect 520920 349757 520980 350106
rect 523368 349890 523428 350106
rect 525952 349890 526012 350106
rect 523358 349830 523428 349890
rect 525934 349830 526012 349890
rect 520917 349756 520983 349757
rect 520917 349692 520918 349756
rect 520982 349692 520983 349756
rect 520917 349691 520983 349692
rect 523358 349077 523418 349830
rect 523355 349076 523421 349077
rect 523355 349012 523356 349076
rect 523420 349012 523421 349076
rect 523355 349011 523421 349012
rect 525934 347717 525994 349830
rect 513419 347716 513485 347717
rect 513419 347652 513420 347716
rect 513484 347652 513485 347716
rect 513419 347651 513485 347652
rect 518387 347716 518453 347717
rect 518387 347652 518388 347716
rect 518452 347652 518453 347716
rect 518387 347651 518453 347652
rect 525931 347716 525997 347717
rect 525931 347652 525932 347716
rect 525996 347652 525997 347716
rect 525931 347651 525997 347652
rect 493363 347172 493429 347173
rect 493363 347108 493364 347172
rect 493428 347108 493429 347172
rect 493363 347107 493429 347108
rect 460611 347036 460677 347037
rect 460611 346972 460612 347036
rect 460676 346972 460677 347036
rect 460611 346971 460677 346972
rect 465947 347036 466013 347037
rect 465947 346972 465948 347036
rect 466012 346972 466013 347036
rect 465947 346971 466013 346972
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 550955 335476 551021 335477
rect 550955 335412 550956 335476
rect 551020 335412 551021 335476
rect 550955 335411 551021 335412
rect 550958 333570 551018 335411
rect 550840 333510 551018 333570
rect 550840 333202 550900 333510
rect 420272 331174 420620 331206
rect 420272 330938 420328 331174
rect 420564 330938 420620 331174
rect 420272 330854 420620 330938
rect 420272 330618 420328 330854
rect 420564 330618 420620 330854
rect 420272 330586 420620 330618
rect 556000 331174 556348 331206
rect 556000 330938 556056 331174
rect 556292 330938 556348 331174
rect 556000 330854 556348 330938
rect 556000 330618 556056 330854
rect 556292 330618 556348 330854
rect 556000 330586 556348 330618
rect 420952 327454 421300 327486
rect 420952 327218 421008 327454
rect 421244 327218 421300 327454
rect 420952 327134 421300 327218
rect 420952 326898 421008 327134
rect 421244 326898 421300 327134
rect 420952 326866 421300 326898
rect 555320 327454 555668 327486
rect 555320 327218 555376 327454
rect 555612 327218 555668 327454
rect 555320 327134 555668 327218
rect 555320 326898 555376 327134
rect 555612 326898 555668 327134
rect 555320 326866 555668 326898
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 420272 295174 420620 295206
rect 420272 294938 420328 295174
rect 420564 294938 420620 295174
rect 420272 294854 420620 294938
rect 420272 294618 420328 294854
rect 420564 294618 420620 294854
rect 420272 294586 420620 294618
rect 556000 295174 556348 295206
rect 556000 294938 556056 295174
rect 556292 294938 556348 295174
rect 556000 294854 556348 294938
rect 556000 294618 556056 294854
rect 556292 294618 556348 294854
rect 556000 294586 556348 294618
rect 420952 291454 421300 291486
rect 420952 291218 421008 291454
rect 421244 291218 421300 291454
rect 420952 291134 421300 291218
rect 420952 290898 421008 291134
rect 421244 290898 421300 291134
rect 420952 290866 421300 290898
rect 555320 291454 555668 291486
rect 555320 291218 555376 291454
rect 555612 291218 555668 291454
rect 555320 291134 555668 291218
rect 555320 290898 555376 291134
rect 555612 290898 555668 291134
rect 555320 290866 555668 290898
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 420272 259174 420620 259206
rect 420272 258938 420328 259174
rect 420564 258938 420620 259174
rect 420272 258854 420620 258938
rect 420272 258618 420328 258854
rect 420564 258618 420620 258854
rect 420272 258586 420620 258618
rect 556000 259174 556348 259206
rect 556000 258938 556056 259174
rect 556292 258938 556348 259174
rect 556000 258854 556348 258938
rect 556000 258618 556056 258854
rect 556292 258618 556348 258854
rect 556000 258586 556348 258618
rect 420952 255454 421300 255486
rect 420952 255218 421008 255454
rect 421244 255218 421300 255454
rect 420952 255134 421300 255218
rect 420952 254898 421008 255134
rect 421244 254898 421300 255134
rect 420952 254866 421300 254898
rect 555320 255454 555668 255486
rect 555320 255218 555376 255454
rect 555612 255218 555668 255454
rect 555320 255134 555668 255218
rect 555320 254898 555376 255134
rect 555612 254898 555668 255134
rect 555320 254866 555668 254898
rect 436056 249930 436116 250106
rect 437144 249930 437204 250106
rect 438232 249930 438292 250106
rect 436056 249870 436202 249930
rect 419766 248370 420010 248430
rect 419950 238645 420010 248370
rect 436142 247077 436202 249870
rect 437062 249870 437204 249930
rect 438166 249870 438292 249930
rect 439592 249930 439652 250106
rect 440544 249930 440604 250106
rect 441768 249930 441828 250106
rect 439592 249870 439698 249930
rect 440544 249870 440618 249930
rect 437062 247349 437122 249870
rect 437059 247348 437125 247349
rect 437059 247284 437060 247348
rect 437124 247284 437125 247348
rect 437059 247283 437125 247284
rect 438166 247077 438226 249870
rect 439638 247077 439698 249870
rect 440558 247077 440618 249870
rect 441662 249870 441828 249930
rect 443128 249930 443188 250106
rect 444216 249930 444276 250106
rect 445440 249930 445500 250106
rect 446528 249930 446588 250106
rect 447616 249930 447676 250106
rect 448296 249930 448356 250106
rect 448704 249930 448764 250106
rect 443128 249870 443194 249930
rect 444216 249870 444298 249930
rect 445440 249870 445586 249930
rect 446528 249870 446690 249930
rect 447616 249870 447794 249930
rect 441662 247077 441722 249870
rect 443134 248301 443194 249870
rect 443131 248300 443197 248301
rect 443131 248236 443132 248300
rect 443196 248236 443197 248300
rect 443131 248235 443197 248236
rect 444238 247077 444298 249870
rect 445526 247077 445586 249870
rect 446630 247077 446690 249870
rect 447734 247077 447794 249870
rect 448286 249870 448356 249930
rect 448654 249870 448764 249930
rect 450064 249930 450124 250106
rect 450744 249930 450804 250106
rect 451288 249930 451348 250106
rect 450064 249870 450186 249930
rect 448286 248301 448346 249870
rect 448654 248301 448714 249870
rect 450126 248301 450186 249870
rect 450678 249870 450804 249930
rect 451046 249870 451348 249930
rect 450678 248301 450738 249870
rect 451046 248430 451106 249870
rect 452376 249658 452436 250106
rect 453464 249658 453524 250106
rect 452334 249598 452436 249658
rect 453438 249598 453524 249658
rect 453600 249658 453660 250106
rect 454552 249658 454612 250106
rect 455912 249658 455972 250106
rect 453600 249598 453682 249658
rect 451046 248370 451290 248430
rect 451230 248301 451290 248370
rect 448283 248300 448349 248301
rect 448283 248236 448284 248300
rect 448348 248236 448349 248300
rect 448283 248235 448349 248236
rect 448651 248300 448717 248301
rect 448651 248236 448652 248300
rect 448716 248236 448717 248300
rect 448651 248235 448717 248236
rect 450123 248300 450189 248301
rect 450123 248236 450124 248300
rect 450188 248236 450189 248300
rect 450123 248235 450189 248236
rect 450675 248300 450741 248301
rect 450675 248236 450676 248300
rect 450740 248236 450741 248300
rect 450675 248235 450741 248236
rect 451227 248300 451293 248301
rect 451227 248236 451228 248300
rect 451292 248236 451293 248300
rect 451227 248235 451293 248236
rect 452334 247077 452394 249598
rect 453438 247077 453498 249598
rect 453622 248301 453682 249598
rect 454542 249598 454612 249658
rect 455830 249598 455972 249658
rect 456048 249658 456108 250106
rect 457000 249658 457060 250106
rect 458088 249658 458148 250106
rect 458496 249658 458556 250106
rect 456048 249598 456258 249658
rect 457000 249598 457178 249658
rect 453619 248300 453685 248301
rect 453619 248236 453620 248300
rect 453684 248236 453685 248300
rect 453619 248235 453685 248236
rect 454542 247077 454602 249598
rect 455830 247621 455890 249598
rect 456198 248301 456258 249598
rect 456195 248300 456261 248301
rect 456195 248236 456196 248300
rect 456260 248236 456261 248300
rect 456195 248235 456261 248236
rect 455827 247620 455893 247621
rect 455827 247556 455828 247620
rect 455892 247556 455893 247620
rect 455827 247555 455893 247556
rect 457118 247349 457178 249598
rect 458038 249598 458148 249658
rect 458406 249598 458556 249658
rect 459448 249658 459508 250106
rect 460672 249658 460732 250106
rect 461080 249661 461140 250106
rect 461760 249930 461820 250106
rect 462848 249930 462908 250106
rect 461718 249870 461820 249930
rect 462822 249870 462908 249930
rect 463528 249930 463588 250106
rect 463936 249930 463996 250106
rect 465296 249930 465356 250106
rect 465976 249930 466036 250106
rect 466384 249930 466444 250106
rect 467608 249930 467668 250106
rect 463528 249870 463618 249930
rect 459448 249598 459570 249658
rect 457115 247348 457181 247349
rect 457115 247284 457116 247348
rect 457180 247284 457181 247348
rect 457115 247283 457181 247284
rect 458038 247077 458098 249598
rect 458406 247757 458466 249598
rect 458403 247756 458469 247757
rect 458403 247692 458404 247756
rect 458468 247692 458469 247756
rect 458403 247691 458469 247692
rect 459510 247349 459570 249598
rect 460614 249598 460732 249658
rect 461077 249660 461143 249661
rect 460614 247621 460674 249598
rect 461077 249596 461078 249660
rect 461142 249596 461143 249660
rect 461077 249595 461143 249596
rect 461718 248029 461778 249870
rect 462822 248301 462882 249870
rect 462819 248300 462885 248301
rect 462819 248236 462820 248300
rect 462884 248236 462885 248300
rect 462819 248235 462885 248236
rect 461715 248028 461781 248029
rect 461715 247964 461716 248028
rect 461780 247964 461781 248028
rect 461715 247963 461781 247964
rect 463558 247893 463618 249870
rect 463926 249870 463996 249930
rect 465214 249870 465356 249930
rect 465950 249870 466036 249930
rect 466318 249870 466444 249930
rect 467606 249870 467668 249930
rect 463926 247893 463986 249870
rect 465214 248029 465274 249870
rect 465211 248028 465277 248029
rect 465211 247964 465212 248028
rect 465276 247964 465277 248028
rect 465211 247963 465277 247964
rect 463555 247892 463621 247893
rect 463555 247828 463556 247892
rect 463620 247828 463621 247892
rect 463555 247827 463621 247828
rect 463923 247892 463989 247893
rect 463923 247828 463924 247892
rect 463988 247828 463989 247892
rect 463923 247827 463989 247828
rect 465950 247757 466010 249870
rect 465947 247756 466013 247757
rect 465947 247692 465948 247756
rect 466012 247692 466013 247756
rect 465947 247691 466013 247692
rect 466318 247621 466378 249870
rect 467606 247757 467666 249870
rect 468288 249797 468348 250106
rect 468696 249930 468756 250106
rect 469784 249930 469844 250106
rect 468696 249870 468770 249930
rect 469784 249870 469874 249930
rect 468285 249796 468351 249797
rect 468285 249732 468286 249796
rect 468350 249732 468351 249796
rect 468285 249731 468351 249732
rect 468710 248301 468770 249870
rect 468707 248300 468773 248301
rect 468707 248236 468708 248300
rect 468772 248236 468773 248300
rect 468707 248235 468773 248236
rect 469814 247893 469874 249870
rect 471008 249661 471068 250106
rect 471144 249930 471204 250106
rect 472232 249930 472292 250106
rect 473320 249930 473380 250106
rect 471144 249870 471346 249930
rect 471005 249660 471071 249661
rect 471005 249596 471006 249660
rect 471070 249596 471071 249660
rect 471005 249595 471071 249596
rect 469811 247892 469877 247893
rect 469811 247828 469812 247892
rect 469876 247828 469877 247892
rect 469811 247827 469877 247828
rect 467603 247756 467669 247757
rect 467603 247692 467604 247756
rect 467668 247692 467669 247756
rect 467603 247691 467669 247692
rect 471286 247621 471346 249870
rect 472206 249870 472292 249930
rect 473310 249870 473380 249930
rect 473592 249930 473652 250106
rect 474408 249930 474468 250106
rect 475768 249930 475828 250106
rect 473592 249870 473738 249930
rect 474408 249870 474474 249930
rect 460611 247620 460677 247621
rect 460611 247556 460612 247620
rect 460676 247556 460677 247620
rect 460611 247555 460677 247556
rect 466315 247620 466381 247621
rect 466315 247556 466316 247620
rect 466380 247556 466381 247620
rect 466315 247555 466381 247556
rect 471283 247620 471349 247621
rect 471283 247556 471284 247620
rect 471348 247556 471349 247620
rect 471283 247555 471349 247556
rect 472206 247349 472266 249870
rect 473310 247349 473370 249870
rect 473678 249389 473738 249870
rect 473675 249388 473741 249389
rect 473675 249324 473676 249388
rect 473740 249324 473741 249388
rect 473675 249323 473741 249324
rect 474414 247893 474474 249870
rect 475702 249870 475828 249930
rect 476040 249930 476100 250106
rect 476992 249930 477052 250106
rect 476040 249870 476130 249930
rect 474411 247892 474477 247893
rect 474411 247828 474412 247892
rect 474476 247828 474477 247892
rect 474411 247827 474477 247828
rect 475702 247485 475762 249870
rect 476070 249525 476130 249870
rect 476990 249870 477052 249930
rect 478080 249930 478140 250106
rect 478488 249930 478548 250106
rect 478080 249870 478154 249930
rect 476067 249524 476133 249525
rect 476067 249460 476068 249524
rect 476132 249460 476133 249524
rect 476067 249459 476133 249460
rect 476990 247485 477050 249870
rect 475699 247484 475765 247485
rect 475699 247420 475700 247484
rect 475764 247420 475765 247484
rect 475699 247419 475765 247420
rect 476987 247484 477053 247485
rect 476987 247420 476988 247484
rect 477052 247420 477053 247484
rect 476987 247419 477053 247420
rect 478094 247349 478154 249870
rect 478462 249870 478548 249930
rect 479168 249930 479228 250106
rect 480936 249930 480996 250106
rect 479168 249870 479258 249930
rect 478462 248165 478522 249870
rect 478459 248164 478525 248165
rect 478459 248100 478460 248164
rect 478524 248100 478525 248164
rect 478459 248099 478525 248100
rect 479198 247757 479258 249870
rect 480854 249870 480996 249930
rect 479195 247756 479261 247757
rect 479195 247692 479196 247756
rect 479260 247692 479261 247756
rect 479195 247691 479261 247692
rect 459507 247348 459573 247349
rect 459507 247284 459508 247348
rect 459572 247284 459573 247348
rect 459507 247283 459573 247284
rect 472203 247348 472269 247349
rect 472203 247284 472204 247348
rect 472268 247284 472269 247348
rect 472203 247283 472269 247284
rect 473307 247348 473373 247349
rect 473307 247284 473308 247348
rect 473372 247284 473373 247348
rect 473307 247283 473373 247284
rect 478091 247348 478157 247349
rect 478091 247284 478092 247348
rect 478156 247284 478157 247348
rect 478091 247283 478157 247284
rect 480854 247077 480914 249870
rect 483520 249661 483580 250106
rect 485968 249797 486028 250106
rect 488280 249797 488340 250106
rect 491000 249797 491060 250106
rect 493448 249930 493508 250106
rect 493366 249870 493508 249930
rect 485965 249796 486031 249797
rect 485965 249732 485966 249796
rect 486030 249732 486031 249796
rect 485965 249731 486031 249732
rect 488277 249796 488343 249797
rect 488277 249732 488278 249796
rect 488342 249732 488343 249796
rect 488277 249731 488343 249732
rect 490997 249796 491063 249797
rect 490997 249732 490998 249796
rect 491062 249732 491063 249796
rect 490997 249731 491063 249732
rect 483517 249660 483583 249661
rect 483517 249596 483518 249660
rect 483582 249596 483583 249660
rect 483517 249595 483583 249596
rect 493366 247077 493426 249870
rect 495896 249797 495956 250106
rect 498480 249797 498540 250106
rect 500928 249797 500988 250106
rect 503512 249797 503572 250106
rect 495893 249796 495959 249797
rect 495893 249732 495894 249796
rect 495958 249732 495959 249796
rect 495893 249731 495959 249732
rect 498477 249796 498543 249797
rect 498477 249732 498478 249796
rect 498542 249732 498543 249796
rect 498477 249731 498543 249732
rect 500925 249796 500991 249797
rect 500925 249732 500926 249796
rect 500990 249732 500991 249796
rect 500925 249731 500991 249732
rect 503509 249796 503575 249797
rect 503509 249732 503510 249796
rect 503574 249732 503575 249796
rect 503509 249731 503575 249732
rect 505960 249661 506020 250106
rect 508544 249661 508604 250106
rect 510992 249930 511052 250106
rect 513440 249930 513500 250106
rect 510992 249870 511090 249930
rect 505957 249660 506023 249661
rect 505957 249596 505958 249660
rect 506022 249596 506023 249660
rect 505957 249595 506023 249596
rect 508541 249660 508607 249661
rect 508541 249596 508542 249660
rect 508606 249596 508607 249660
rect 508541 249595 508607 249596
rect 511030 247077 511090 249870
rect 513422 249870 513500 249930
rect 513422 247077 513482 249870
rect 515888 249661 515948 250106
rect 518472 249930 518532 250106
rect 518390 249870 518532 249930
rect 515885 249660 515951 249661
rect 515885 249596 515886 249660
rect 515950 249596 515951 249660
rect 515885 249595 515951 249596
rect 518390 247213 518450 249870
rect 520920 249661 520980 250106
rect 523368 249930 523428 250106
rect 525952 249930 526012 250106
rect 523358 249870 523428 249930
rect 525934 249870 526012 249930
rect 520917 249660 520983 249661
rect 520917 249596 520918 249660
rect 520982 249596 520983 249660
rect 520917 249595 520983 249596
rect 518387 247212 518453 247213
rect 518387 247148 518388 247212
rect 518452 247148 518453 247212
rect 518387 247147 518453 247148
rect 523358 247077 523418 249870
rect 525934 247077 525994 249870
rect 436139 247076 436205 247077
rect 436139 247012 436140 247076
rect 436204 247012 436205 247076
rect 436139 247011 436205 247012
rect 438163 247076 438229 247077
rect 438163 247012 438164 247076
rect 438228 247012 438229 247076
rect 438163 247011 438229 247012
rect 439635 247076 439701 247077
rect 439635 247012 439636 247076
rect 439700 247012 439701 247076
rect 439635 247011 439701 247012
rect 440555 247076 440621 247077
rect 440555 247012 440556 247076
rect 440620 247012 440621 247076
rect 440555 247011 440621 247012
rect 441659 247076 441725 247077
rect 441659 247012 441660 247076
rect 441724 247012 441725 247076
rect 441659 247011 441725 247012
rect 444235 247076 444301 247077
rect 444235 247012 444236 247076
rect 444300 247012 444301 247076
rect 444235 247011 444301 247012
rect 445523 247076 445589 247077
rect 445523 247012 445524 247076
rect 445588 247012 445589 247076
rect 445523 247011 445589 247012
rect 446627 247076 446693 247077
rect 446627 247012 446628 247076
rect 446692 247012 446693 247076
rect 446627 247011 446693 247012
rect 447731 247076 447797 247077
rect 447731 247012 447732 247076
rect 447796 247012 447797 247076
rect 447731 247011 447797 247012
rect 452331 247076 452397 247077
rect 452331 247012 452332 247076
rect 452396 247012 452397 247076
rect 452331 247011 452397 247012
rect 453435 247076 453501 247077
rect 453435 247012 453436 247076
rect 453500 247012 453501 247076
rect 453435 247011 453501 247012
rect 454539 247076 454605 247077
rect 454539 247012 454540 247076
rect 454604 247012 454605 247076
rect 454539 247011 454605 247012
rect 458035 247076 458101 247077
rect 458035 247012 458036 247076
rect 458100 247012 458101 247076
rect 458035 247011 458101 247012
rect 480851 247076 480917 247077
rect 480851 247012 480852 247076
rect 480916 247012 480917 247076
rect 480851 247011 480917 247012
rect 493363 247076 493429 247077
rect 493363 247012 493364 247076
rect 493428 247012 493429 247076
rect 493363 247011 493429 247012
rect 511027 247076 511093 247077
rect 511027 247012 511028 247076
rect 511092 247012 511093 247076
rect 511027 247011 511093 247012
rect 513419 247076 513485 247077
rect 513419 247012 513420 247076
rect 513484 247012 513485 247076
rect 513419 247011 513485 247012
rect 523355 247076 523421 247077
rect 523355 247012 523356 247076
rect 523420 247012 523421 247076
rect 523355 247011 523421 247012
rect 525931 247076 525997 247077
rect 525931 247012 525932 247076
rect 525996 247012 525997 247076
rect 525931 247011 525997 247012
rect 419947 238644 420013 238645
rect 419947 238580 419948 238644
rect 420012 238580 420013 238644
rect 419947 238579 420013 238580
rect 419579 235788 419645 235789
rect 419579 235724 419580 235788
rect 419644 235724 419645 235788
rect 419579 235723 419645 235724
rect 419582 234970 419642 235723
rect 419398 234910 419642 234970
rect 419398 147253 419458 234910
rect 419950 148341 420010 238579
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 550771 235108 550837 235109
rect 550771 235044 550772 235108
rect 550836 235044 550837 235108
rect 550771 235043 550837 235044
rect 550774 233610 550834 235043
rect 550774 233550 550900 233610
rect 550840 233240 550900 233550
rect 420272 223174 420620 223206
rect 420272 222938 420328 223174
rect 420564 222938 420620 223174
rect 420272 222854 420620 222938
rect 420272 222618 420328 222854
rect 420564 222618 420620 222854
rect 420272 222586 420620 222618
rect 556000 223174 556348 223206
rect 556000 222938 556056 223174
rect 556292 222938 556348 223174
rect 556000 222854 556348 222938
rect 556000 222618 556056 222854
rect 556292 222618 556348 222854
rect 556000 222586 556348 222618
rect 420952 219454 421300 219486
rect 420952 219218 421008 219454
rect 421244 219218 421300 219454
rect 420952 219134 421300 219218
rect 420952 218898 421008 219134
rect 421244 218898 421300 219134
rect 420952 218866 421300 218898
rect 555320 219454 555668 219486
rect 555320 219218 555376 219454
rect 555612 219218 555668 219454
rect 555320 219134 555668 219218
rect 555320 218898 555376 219134
rect 555612 218898 555668 219134
rect 555320 218866 555668 218898
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 420272 187174 420620 187206
rect 420272 186938 420328 187174
rect 420564 186938 420620 187174
rect 420272 186854 420620 186938
rect 420272 186618 420328 186854
rect 420564 186618 420620 186854
rect 420272 186586 420620 186618
rect 556000 187174 556348 187206
rect 556000 186938 556056 187174
rect 556292 186938 556348 187174
rect 556000 186854 556348 186938
rect 556000 186618 556056 186854
rect 556292 186618 556348 186854
rect 556000 186586 556348 186618
rect 420952 183454 421300 183486
rect 420952 183218 421008 183454
rect 421244 183218 421300 183454
rect 420952 183134 421300 183218
rect 420952 182898 421008 183134
rect 421244 182898 421300 183134
rect 420952 182866 421300 182898
rect 555320 183454 555668 183486
rect 555320 183218 555376 183454
rect 555612 183218 555668 183454
rect 555320 183134 555668 183218
rect 555320 182898 555376 183134
rect 555612 182898 555668 183134
rect 555320 182866 555668 182898
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 420272 151174 420620 151206
rect 420272 150938 420328 151174
rect 420564 150938 420620 151174
rect 420272 150854 420620 150938
rect 420272 150618 420328 150854
rect 420564 150618 420620 150854
rect 420272 150586 420620 150618
rect 556000 151174 556348 151206
rect 556000 150938 556056 151174
rect 556292 150938 556348 151174
rect 556000 150854 556348 150938
rect 556000 150618 556056 150854
rect 556292 150618 556348 150854
rect 556000 150586 556348 150618
rect 436056 149290 436116 150106
rect 437144 149290 437204 150106
rect 438232 149290 438292 150106
rect 436056 149230 436202 149290
rect 419947 148340 420013 148341
rect 419947 148276 419948 148340
rect 420012 148276 420013 148340
rect 419947 148275 420013 148276
rect 419395 147252 419461 147253
rect 419395 147188 419396 147252
rect 419460 147188 419461 147252
rect 419395 147187 419461 147188
rect 419211 146844 419277 146845
rect 419211 146780 419212 146844
rect 419276 146780 419277 146844
rect 419211 146779 419277 146780
rect 418659 49196 418725 49197
rect 418659 49132 418660 49196
rect 418724 49132 418725 49196
rect 418659 49131 418725 49132
rect 419214 47565 419274 146779
rect 419398 48109 419458 147187
rect 419950 49061 420010 148275
rect 436142 147661 436202 149230
rect 437062 149230 437204 149290
rect 438166 149230 438292 149290
rect 439592 149290 439652 150106
rect 440544 149701 440604 150106
rect 440541 149700 440607 149701
rect 440541 149636 440542 149700
rect 440606 149636 440607 149700
rect 440541 149635 440607 149636
rect 441768 149565 441828 150106
rect 441765 149564 441831 149565
rect 441765 149500 441766 149564
rect 441830 149500 441831 149564
rect 441765 149499 441831 149500
rect 443128 149290 443188 150106
rect 444216 149290 444276 150106
rect 445440 149290 445500 150106
rect 446528 149290 446588 150106
rect 447616 149290 447676 150106
rect 448296 149290 448356 150106
rect 448704 149290 448764 150106
rect 439592 149230 439698 149290
rect 443128 149230 443194 149290
rect 444216 149230 444298 149290
rect 437062 147661 437122 149230
rect 438166 147690 438226 149230
rect 437982 147661 438226 147690
rect 439638 147661 439698 149230
rect 443134 147661 443194 149230
rect 444238 147661 444298 149230
rect 445342 149230 445500 149290
rect 446446 149230 446588 149290
rect 447550 149230 447676 149290
rect 448286 149230 448356 149290
rect 448654 149230 448764 149290
rect 450064 149290 450124 150106
rect 450744 149290 450804 150106
rect 451288 149290 451348 150106
rect 452376 149290 452436 150106
rect 453464 149290 453524 150106
rect 450064 149230 450186 149290
rect 445342 147661 445402 149230
rect 446446 147661 446506 149230
rect 447550 147690 447610 149230
rect 447366 147661 447610 147690
rect 448286 147661 448346 149230
rect 448654 147661 448714 149230
rect 450126 147661 450186 149230
rect 450678 149230 450804 149290
rect 451230 149230 451348 149290
rect 452334 149230 452436 149290
rect 453438 149230 453524 149290
rect 453600 149290 453660 150106
rect 454552 149290 454612 150106
rect 455912 149565 455972 150106
rect 455909 149564 455975 149565
rect 455909 149500 455910 149564
rect 455974 149500 455975 149564
rect 455909 149499 455975 149500
rect 456048 149290 456108 150106
rect 457000 149290 457060 150106
rect 458088 149837 458148 150106
rect 458085 149836 458151 149837
rect 458085 149772 458086 149836
rect 458150 149772 458151 149836
rect 458085 149771 458151 149772
rect 458496 149290 458556 150106
rect 453600 149230 453682 149290
rect 450678 147661 450738 149230
rect 451230 147661 451290 149230
rect 452334 147661 452394 149230
rect 453438 147661 453498 149230
rect 453622 147661 453682 149230
rect 454542 149230 454612 149290
rect 456014 149230 456108 149290
rect 456934 149230 457060 149290
rect 458406 149230 458556 149290
rect 459448 149290 459508 150106
rect 460672 149290 460732 150106
rect 461080 149565 461140 150106
rect 461077 149564 461143 149565
rect 461077 149500 461078 149564
rect 461142 149500 461143 149564
rect 461077 149499 461143 149500
rect 461760 149290 461820 150106
rect 462848 149290 462908 150106
rect 463528 149565 463588 150106
rect 463525 149564 463591 149565
rect 463525 149500 463526 149564
rect 463590 149500 463591 149564
rect 463525 149499 463591 149500
rect 463936 149290 463996 150106
rect 465296 149290 465356 150106
rect 465976 149565 466036 150106
rect 465973 149564 466039 149565
rect 465973 149500 465974 149564
rect 466038 149500 466039 149564
rect 465973 149499 466039 149500
rect 466384 149290 466444 150106
rect 467608 149290 467668 150106
rect 468288 149565 468348 150106
rect 468285 149564 468351 149565
rect 468285 149500 468286 149564
rect 468350 149500 468351 149564
rect 468285 149499 468351 149500
rect 459448 149230 459570 149290
rect 454542 147661 454602 149230
rect 456014 147661 456074 149230
rect 436139 147660 436205 147661
rect 436139 147596 436140 147660
rect 436204 147596 436205 147660
rect 436139 147595 436205 147596
rect 437059 147660 437125 147661
rect 437059 147596 437060 147660
rect 437124 147596 437125 147660
rect 437059 147595 437125 147596
rect 437979 147660 438226 147661
rect 437979 147596 437980 147660
rect 438044 147630 438226 147660
rect 439635 147660 439701 147661
rect 438044 147596 438045 147630
rect 437979 147595 438045 147596
rect 439635 147596 439636 147660
rect 439700 147596 439701 147660
rect 439635 147595 439701 147596
rect 443131 147660 443197 147661
rect 443131 147596 443132 147660
rect 443196 147596 443197 147660
rect 443131 147595 443197 147596
rect 444235 147660 444301 147661
rect 444235 147596 444236 147660
rect 444300 147596 444301 147660
rect 444235 147595 444301 147596
rect 445339 147660 445405 147661
rect 445339 147596 445340 147660
rect 445404 147596 445405 147660
rect 445339 147595 445405 147596
rect 446443 147660 446509 147661
rect 446443 147596 446444 147660
rect 446508 147596 446509 147660
rect 446443 147595 446509 147596
rect 447363 147660 447610 147661
rect 447363 147596 447364 147660
rect 447428 147630 447610 147660
rect 448283 147660 448349 147661
rect 447428 147596 447429 147630
rect 447363 147595 447429 147596
rect 448283 147596 448284 147660
rect 448348 147596 448349 147660
rect 448283 147595 448349 147596
rect 448651 147660 448717 147661
rect 448651 147596 448652 147660
rect 448716 147596 448717 147660
rect 448651 147595 448717 147596
rect 450123 147660 450189 147661
rect 450123 147596 450124 147660
rect 450188 147596 450189 147660
rect 450123 147595 450189 147596
rect 450675 147660 450741 147661
rect 450675 147596 450676 147660
rect 450740 147596 450741 147660
rect 450675 147595 450741 147596
rect 451227 147660 451293 147661
rect 451227 147596 451228 147660
rect 451292 147596 451293 147660
rect 451227 147595 451293 147596
rect 452331 147660 452397 147661
rect 452331 147596 452332 147660
rect 452396 147596 452397 147660
rect 452331 147595 452397 147596
rect 453435 147660 453501 147661
rect 453435 147596 453436 147660
rect 453500 147596 453501 147660
rect 453435 147595 453501 147596
rect 453619 147660 453685 147661
rect 453619 147596 453620 147660
rect 453684 147596 453685 147660
rect 453619 147595 453685 147596
rect 454539 147660 454605 147661
rect 454539 147596 454540 147660
rect 454604 147596 454605 147660
rect 454539 147595 454605 147596
rect 456011 147660 456077 147661
rect 456011 147596 456012 147660
rect 456076 147596 456077 147660
rect 456011 147595 456077 147596
rect 456934 147117 456994 149230
rect 458406 147661 458466 149230
rect 459510 148749 459570 149230
rect 460614 149230 460732 149290
rect 461718 149230 461820 149290
rect 462822 149230 462908 149290
rect 463926 149230 463996 149290
rect 465214 149230 465356 149290
rect 466318 149230 466444 149290
rect 467606 149230 467668 149290
rect 468696 149290 468756 150106
rect 469784 149290 469844 150106
rect 471008 149565 471068 150106
rect 471005 149564 471071 149565
rect 471005 149500 471006 149564
rect 471070 149500 471071 149564
rect 471005 149499 471071 149500
rect 471144 149290 471204 150106
rect 472232 149290 472292 150106
rect 473320 149290 473380 150106
rect 473592 149290 473652 150106
rect 468696 149230 468770 149290
rect 469784 149230 469874 149290
rect 459507 148748 459573 148749
rect 459507 148684 459508 148748
rect 459572 148684 459573 148748
rect 459507 148683 459573 148684
rect 458403 147660 458469 147661
rect 458403 147596 458404 147660
rect 458468 147596 458469 147660
rect 458403 147595 458469 147596
rect 456931 147116 456997 147117
rect 456931 147052 456932 147116
rect 456996 147052 456997 147116
rect 456931 147051 456997 147052
rect 456934 146845 456994 147051
rect 460614 146981 460674 149230
rect 461718 147661 461778 149230
rect 462822 147661 462882 149230
rect 463926 147661 463986 149230
rect 465214 147661 465274 149230
rect 466318 147661 466378 149230
rect 467606 147661 467666 149230
rect 468710 147661 468770 149230
rect 469814 147661 469874 149230
rect 471102 149230 471204 149290
rect 472206 149230 472292 149290
rect 473310 149230 473380 149290
rect 473494 149230 473652 149290
rect 474408 149290 474468 150106
rect 475768 149290 475828 150106
rect 476040 149834 476100 150106
rect 476992 149834 477052 150106
rect 476040 149774 476130 149834
rect 474408 149230 474474 149290
rect 471102 147661 471162 149230
rect 472206 147661 472266 149230
rect 473310 147661 473370 149230
rect 461715 147660 461781 147661
rect 461715 147596 461716 147660
rect 461780 147596 461781 147660
rect 461715 147595 461781 147596
rect 462819 147660 462885 147661
rect 462819 147596 462820 147660
rect 462884 147596 462885 147660
rect 462819 147595 462885 147596
rect 463923 147660 463989 147661
rect 463923 147596 463924 147660
rect 463988 147596 463989 147660
rect 463923 147595 463989 147596
rect 465211 147660 465277 147661
rect 465211 147596 465212 147660
rect 465276 147596 465277 147660
rect 465211 147595 465277 147596
rect 466315 147660 466381 147661
rect 466315 147596 466316 147660
rect 466380 147596 466381 147660
rect 466315 147595 466381 147596
rect 467603 147660 467669 147661
rect 467603 147596 467604 147660
rect 467668 147596 467669 147660
rect 467603 147595 467669 147596
rect 468707 147660 468773 147661
rect 468707 147596 468708 147660
rect 468772 147596 468773 147660
rect 468707 147595 468773 147596
rect 469811 147660 469877 147661
rect 469811 147596 469812 147660
rect 469876 147596 469877 147660
rect 469811 147595 469877 147596
rect 471099 147660 471165 147661
rect 471099 147596 471100 147660
rect 471164 147596 471165 147660
rect 471099 147595 471165 147596
rect 472203 147660 472269 147661
rect 472203 147596 472204 147660
rect 472268 147596 472269 147660
rect 472203 147595 472269 147596
rect 473307 147660 473373 147661
rect 473307 147596 473308 147660
rect 473372 147596 473373 147660
rect 473307 147595 473373 147596
rect 473494 147253 473554 149230
rect 474414 147661 474474 149230
rect 475702 149230 475828 149290
rect 475702 147690 475762 149230
rect 476070 149157 476130 149774
rect 476990 149774 477052 149834
rect 478080 149834 478140 150106
rect 478488 149837 478548 150106
rect 478485 149836 478551 149837
rect 478080 149774 478154 149834
rect 476067 149156 476133 149157
rect 476067 149092 476068 149156
rect 476132 149092 476133 149156
rect 476067 149091 476133 149092
rect 474411 147660 474477 147661
rect 474411 147596 474412 147660
rect 474476 147596 474477 147660
rect 474411 147595 474477 147596
rect 475518 147630 475762 147690
rect 476990 147661 477050 149774
rect 478094 147661 478154 149774
rect 478485 149772 478486 149836
rect 478550 149772 478551 149836
rect 479168 149834 479228 150106
rect 480936 149837 480996 150106
rect 483520 149837 483580 150106
rect 485968 149837 486028 150106
rect 480933 149836 480999 149837
rect 479168 149774 479258 149834
rect 478485 149771 478551 149772
rect 476987 147660 477053 147661
rect 473491 147252 473557 147253
rect 473491 147188 473492 147252
rect 473556 147188 473557 147252
rect 473491 147187 473557 147188
rect 460611 146980 460677 146981
rect 460611 146916 460612 146980
rect 460676 146916 460677 146980
rect 460611 146915 460677 146916
rect 475518 146845 475578 147630
rect 476987 147596 476988 147660
rect 477052 147596 477053 147660
rect 476987 147595 477053 147596
rect 478091 147660 478157 147661
rect 478091 147596 478092 147660
rect 478156 147596 478157 147660
rect 478091 147595 478157 147596
rect 479198 147117 479258 149774
rect 480933 149772 480934 149836
rect 480998 149772 480999 149836
rect 480933 149771 480999 149772
rect 483517 149836 483583 149837
rect 483517 149772 483518 149836
rect 483582 149772 483583 149836
rect 483517 149771 483583 149772
rect 485965 149836 486031 149837
rect 485965 149772 485966 149836
rect 486030 149772 486031 149836
rect 485965 149771 486031 149772
rect 488280 149701 488340 150106
rect 491000 149701 491060 150106
rect 488277 149700 488343 149701
rect 488277 149636 488278 149700
rect 488342 149636 488343 149700
rect 488277 149635 488343 149636
rect 490997 149700 491063 149701
rect 490997 149636 490998 149700
rect 491062 149636 491063 149700
rect 490997 149635 491063 149636
rect 493448 149290 493508 150106
rect 495896 149701 495956 150106
rect 495893 149700 495959 149701
rect 495893 149636 495894 149700
rect 495958 149636 495959 149700
rect 495893 149635 495959 149636
rect 493366 149230 493508 149290
rect 498480 149290 498540 150106
rect 500928 149290 500988 150106
rect 503512 149701 503572 150106
rect 503509 149700 503575 149701
rect 503509 149636 503510 149700
rect 503574 149636 503575 149700
rect 503509 149635 503575 149636
rect 505960 149565 506020 150106
rect 508544 149565 508604 150106
rect 510992 149565 511052 150106
rect 505957 149564 506023 149565
rect 505957 149500 505958 149564
rect 506022 149500 506023 149564
rect 505957 149499 506023 149500
rect 508541 149564 508607 149565
rect 508541 149500 508542 149564
rect 508606 149500 508607 149564
rect 508541 149499 508607 149500
rect 510989 149564 511055 149565
rect 510989 149500 510990 149564
rect 511054 149500 511055 149564
rect 510989 149499 511055 149500
rect 513440 149290 513500 150106
rect 515888 149565 515948 150106
rect 518472 149565 518532 150106
rect 515885 149564 515951 149565
rect 515885 149500 515886 149564
rect 515950 149500 515951 149564
rect 515885 149499 515951 149500
rect 518469 149564 518535 149565
rect 518469 149500 518470 149564
rect 518534 149500 518535 149564
rect 520920 149562 520980 150106
rect 523368 149562 523428 150106
rect 525952 149562 526012 150106
rect 520920 149502 521026 149562
rect 518469 149499 518535 149500
rect 498480 149230 498578 149290
rect 493366 147389 493426 149230
rect 493363 147388 493429 147389
rect 493363 147324 493364 147388
rect 493428 147324 493429 147388
rect 493363 147323 493429 147324
rect 479195 147116 479261 147117
rect 479195 147052 479196 147116
rect 479260 147052 479261 147116
rect 479195 147051 479261 147052
rect 456931 146844 456997 146845
rect 456931 146780 456932 146844
rect 456996 146780 456997 146844
rect 456931 146779 456997 146780
rect 475515 146844 475581 146845
rect 475515 146780 475516 146844
rect 475580 146780 475581 146844
rect 475515 146779 475581 146780
rect 498518 146573 498578 149230
rect 500910 149230 500988 149290
rect 513422 149230 513500 149290
rect 500910 147525 500970 149230
rect 513422 149021 513482 149230
rect 520966 149021 521026 149502
rect 523358 149502 523428 149562
rect 525934 149502 526012 149562
rect 523358 149021 523418 149502
rect 525934 149021 525994 149502
rect 513419 149020 513485 149021
rect 513419 148956 513420 149020
rect 513484 148956 513485 149020
rect 513419 148955 513485 148956
rect 520963 149020 521029 149021
rect 520963 148956 520964 149020
rect 521028 148956 521029 149020
rect 520963 148955 521029 148956
rect 523355 149020 523421 149021
rect 523355 148956 523356 149020
rect 523420 148956 523421 149020
rect 523355 148955 523421 148956
rect 525931 149020 525997 149021
rect 525931 148956 525932 149020
rect 525996 148956 525997 149020
rect 525931 148955 525997 148956
rect 500907 147524 500973 147525
rect 500907 147460 500908 147524
rect 500972 147460 500973 147524
rect 500907 147459 500973 147460
rect 498515 146572 498581 146573
rect 498515 146508 498516 146572
rect 498580 146508 498581 146572
rect 498515 146507 498581 146508
rect 551507 136508 551573 136509
rect 551507 136444 551508 136508
rect 551572 136444 551573 136508
rect 551507 136443 551573 136444
rect 551510 133310 551570 136443
rect 550870 133250 551570 133310
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 420272 115174 420620 115206
rect 420272 114938 420328 115174
rect 420564 114938 420620 115174
rect 420272 114854 420620 114938
rect 420272 114618 420328 114854
rect 420564 114618 420620 114854
rect 420272 114586 420620 114618
rect 556000 115174 556348 115206
rect 556000 114938 556056 115174
rect 556292 114938 556348 115174
rect 556000 114854 556348 114938
rect 556000 114618 556056 114854
rect 556292 114618 556348 114854
rect 556000 114586 556348 114618
rect 420952 111454 421300 111486
rect 420952 111218 421008 111454
rect 421244 111218 421300 111454
rect 420952 111134 421300 111218
rect 420952 110898 421008 111134
rect 421244 110898 421300 111134
rect 420952 110866 421300 110898
rect 555320 111454 555668 111486
rect 555320 111218 555376 111454
rect 555612 111218 555668 111454
rect 555320 111134 555668 111218
rect 555320 110898 555376 111134
rect 555612 110898 555668 111134
rect 555320 110866 555668 110898
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 420272 79174 420620 79206
rect 420272 78938 420328 79174
rect 420564 78938 420620 79174
rect 420272 78854 420620 78938
rect 420272 78618 420328 78854
rect 420564 78618 420620 78854
rect 420272 78586 420620 78618
rect 556000 79174 556348 79206
rect 556000 78938 556056 79174
rect 556292 78938 556348 79174
rect 556000 78854 556348 78938
rect 556000 78618 556056 78854
rect 556292 78618 556348 78854
rect 556000 78586 556348 78618
rect 420952 75454 421300 75486
rect 420952 75218 421008 75454
rect 421244 75218 421300 75454
rect 420952 75134 421300 75218
rect 420952 74898 421008 75134
rect 421244 74898 421300 75134
rect 420952 74866 421300 74898
rect 555320 75454 555668 75486
rect 555320 75218 555376 75454
rect 555612 75218 555668 75454
rect 555320 75134 555668 75218
rect 555320 74898 555376 75134
rect 555612 74898 555668 75134
rect 555320 74866 555668 74898
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 436056 50010 436116 50106
rect 437144 50010 437204 50106
rect 438232 50010 438292 50106
rect 436056 49950 436202 50010
rect 419947 49060 420013 49061
rect 419947 48996 419948 49060
rect 420012 48996 420013 49060
rect 419947 48995 420013 48996
rect 436142 48245 436202 49950
rect 437062 49950 437204 50010
rect 438166 49950 438292 50010
rect 439592 50010 439652 50106
rect 440544 50010 440604 50106
rect 441768 50010 441828 50106
rect 443128 50010 443188 50106
rect 444216 50010 444276 50106
rect 445440 50010 445500 50106
rect 446528 50010 446588 50106
rect 447616 50010 447676 50106
rect 448296 50010 448356 50106
rect 448704 50010 448764 50106
rect 439592 49950 439698 50010
rect 440544 49950 440618 50010
rect 441768 49950 442090 50010
rect 443128 49950 443194 50010
rect 444216 49950 444298 50010
rect 437062 48245 437122 49950
rect 438166 48245 438226 49950
rect 439638 48245 439698 49950
rect 436139 48244 436205 48245
rect 436139 48180 436140 48244
rect 436204 48180 436205 48244
rect 436139 48179 436205 48180
rect 437059 48244 437125 48245
rect 437059 48180 437060 48244
rect 437124 48180 437125 48244
rect 437059 48179 437125 48180
rect 438163 48244 438229 48245
rect 438163 48180 438164 48244
rect 438228 48180 438229 48244
rect 438163 48179 438229 48180
rect 439635 48244 439701 48245
rect 439635 48180 439636 48244
rect 439700 48180 439701 48244
rect 439635 48179 439701 48180
rect 440558 48109 440618 49950
rect 419395 48108 419461 48109
rect 419395 48044 419396 48108
rect 419460 48044 419461 48108
rect 440555 48108 440621 48109
rect 419395 48043 419461 48044
rect 419211 47564 419277 47565
rect 419211 47500 419212 47564
rect 419276 47500 419277 47564
rect 419211 47499 419277 47500
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 25774 420734 48064
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 29494 424454 48064
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 39454 434414 48064
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 43174 438134 48064
rect 440555 48044 440556 48108
rect 440620 48044 440621 48108
rect 440555 48043 440621 48044
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 46894 441854 47940
rect 442030 47429 442090 49950
rect 443134 48245 443194 49950
rect 444238 48245 444298 49950
rect 445342 49950 445500 50010
rect 446446 49950 446588 50010
rect 447550 49950 447676 50010
rect 448286 49950 448356 50010
rect 448654 49950 448764 50010
rect 450064 50010 450124 50106
rect 450744 50010 450804 50106
rect 451288 50010 451348 50106
rect 452376 50010 452436 50106
rect 453464 50010 453524 50106
rect 450064 49950 450186 50010
rect 443131 48244 443197 48245
rect 443131 48180 443132 48244
rect 443196 48180 443197 48244
rect 443131 48179 443197 48180
rect 444235 48244 444301 48245
rect 444235 48180 444236 48244
rect 444300 48180 444301 48244
rect 444235 48179 444301 48180
rect 445342 48109 445402 49950
rect 446446 48109 446506 49950
rect 445339 48108 445405 48109
rect 445339 48044 445340 48108
rect 445404 48044 445405 48108
rect 445339 48043 445405 48044
rect 446443 48108 446509 48109
rect 446443 48044 446444 48108
rect 446508 48044 446509 48108
rect 446443 48043 446509 48044
rect 442027 47428 442093 47429
rect 442027 47364 442028 47428
rect 442092 47364 442093 47428
rect 442027 47363 442093 47364
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 47940
rect 447550 47565 447610 49950
rect 448286 48245 448346 49950
rect 448283 48244 448349 48245
rect 448283 48180 448284 48244
rect 448348 48180 448349 48244
rect 448283 48179 448349 48180
rect 448654 48109 448714 49950
rect 448651 48108 448717 48109
rect 448651 48044 448652 48108
rect 448716 48044 448717 48108
rect 448651 48043 448717 48044
rect 447547 47564 447613 47565
rect 447547 47500 447548 47564
rect 447612 47500 447613 47564
rect 447547 47499 447613 47500
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 47940
rect 450126 47429 450186 49950
rect 450678 49950 450804 50010
rect 451046 49950 451348 50010
rect 452334 49950 452436 50010
rect 453438 49950 453524 50010
rect 453600 50010 453660 50106
rect 454552 50010 454612 50106
rect 455912 50010 455972 50106
rect 453600 49950 453682 50010
rect 450678 48245 450738 49950
rect 450675 48244 450741 48245
rect 450675 48180 450676 48244
rect 450740 48180 450741 48244
rect 450675 48179 450741 48180
rect 450123 47428 450189 47429
rect 450123 47364 450124 47428
rect 450188 47364 450189 47428
rect 450123 47363 450189 47364
rect 451046 47290 451106 49950
rect 452334 48109 452394 49950
rect 453438 48109 453498 49950
rect 453622 48245 453682 49950
rect 454542 49950 454612 50010
rect 455646 49950 455972 50010
rect 454542 48245 454602 49950
rect 455646 48245 455706 49950
rect 456048 49330 456108 50106
rect 457000 49877 457060 50106
rect 458088 49877 458148 50106
rect 458496 50010 458556 50106
rect 458406 49950 458556 50010
rect 459448 50010 459508 50106
rect 460672 50010 460732 50106
rect 461080 50010 461140 50106
rect 461760 50010 461820 50106
rect 462848 50010 462908 50106
rect 459448 49950 459570 50010
rect 456997 49876 457063 49877
rect 456997 49812 456998 49876
rect 457062 49812 457063 49876
rect 456997 49811 457063 49812
rect 458085 49876 458151 49877
rect 458085 49812 458086 49876
rect 458150 49812 458151 49876
rect 458085 49811 458151 49812
rect 455830 49270 456108 49330
rect 453619 48244 453685 48245
rect 453619 48180 453620 48244
rect 453684 48180 453685 48244
rect 453619 48179 453685 48180
rect 454539 48244 454605 48245
rect 454539 48180 454540 48244
rect 454604 48180 454605 48244
rect 454539 48179 454605 48180
rect 455643 48244 455709 48245
rect 455643 48180 455644 48244
rect 455708 48180 455709 48244
rect 455643 48179 455709 48180
rect 452331 48108 452397 48109
rect 452331 48044 452332 48108
rect 452396 48044 452397 48108
rect 452331 48043 452397 48044
rect 453435 48108 453501 48109
rect 453435 48044 453436 48108
rect 453500 48044 453501 48108
rect 453435 48043 453501 48044
rect 451227 47428 451293 47429
rect 451227 47364 451228 47428
rect 451292 47364 451293 47428
rect 451227 47363 451293 47364
rect 451230 47290 451290 47363
rect 451046 47230 451290 47290
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 47940
rect 455830 47701 455890 49270
rect 458406 48245 458466 49950
rect 459510 49061 459570 49950
rect 460614 49950 460732 50010
rect 460982 49950 461140 50010
rect 461718 49950 461820 50010
rect 462822 49950 462908 50010
rect 463528 50010 463588 50106
rect 463936 50010 463996 50106
rect 465296 50010 465356 50106
rect 465976 50010 466036 50106
rect 466384 50010 466444 50106
rect 467608 50010 467668 50106
rect 463528 49950 463618 50010
rect 459507 49060 459573 49061
rect 459507 48996 459508 49060
rect 459572 48996 459573 49060
rect 459507 48995 459573 48996
rect 458403 48244 458469 48245
rect 458403 48180 458404 48244
rect 458468 48180 458469 48244
rect 458403 48179 458469 48180
rect 455827 47700 455893 47701
rect 455827 47636 455828 47700
rect 455892 47636 455893 47700
rect 455827 47635 455893 47636
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 25774 456734 47940
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 48064
rect 460614 47701 460674 49950
rect 460982 49197 461042 49950
rect 460979 49196 461045 49197
rect 460979 49132 460980 49196
rect 461044 49132 461045 49196
rect 460979 49131 461045 49132
rect 461718 48245 461778 49950
rect 462822 48245 462882 49950
rect 463558 48245 463618 49950
rect 463926 49950 463996 50010
rect 465214 49950 465356 50010
rect 465950 49950 466036 50010
rect 466318 49950 466444 50010
rect 467606 49950 467668 50010
rect 468288 50010 468348 50106
rect 468696 50010 468756 50106
rect 469784 50010 469844 50106
rect 468288 49950 468402 50010
rect 468696 49950 468770 50010
rect 469784 49950 469874 50010
rect 463926 48245 463986 49950
rect 465214 48245 465274 49950
rect 465950 48245 466010 49950
rect 466318 48245 466378 49950
rect 467606 48245 467666 49950
rect 468342 48245 468402 49950
rect 468710 48245 468770 49950
rect 469814 48245 469874 49950
rect 471008 49330 471068 50106
rect 471144 50010 471204 50106
rect 472232 50010 472292 50106
rect 471144 49950 471346 50010
rect 470918 49270 471068 49330
rect 470918 48245 470978 49270
rect 471286 48245 471346 49950
rect 472206 49950 472292 50010
rect 472206 48245 472266 49950
rect 473320 49741 473380 50106
rect 473592 50010 473652 50106
rect 473494 49950 473652 50010
rect 474408 50010 474468 50106
rect 475768 50010 475828 50106
rect 474408 49950 474474 50010
rect 473317 49740 473383 49741
rect 473317 49676 473318 49740
rect 473382 49676 473383 49740
rect 473317 49675 473383 49676
rect 473494 49330 473554 49950
rect 473310 49270 473554 49330
rect 461715 48244 461781 48245
rect 461715 48180 461716 48244
rect 461780 48180 461781 48244
rect 461715 48179 461781 48180
rect 462819 48244 462885 48245
rect 462819 48180 462820 48244
rect 462884 48180 462885 48244
rect 462819 48179 462885 48180
rect 463555 48244 463621 48245
rect 463555 48180 463556 48244
rect 463620 48180 463621 48244
rect 463555 48179 463621 48180
rect 463923 48244 463989 48245
rect 463923 48180 463924 48244
rect 463988 48180 463989 48244
rect 463923 48179 463989 48180
rect 465211 48244 465277 48245
rect 465211 48180 465212 48244
rect 465276 48180 465277 48244
rect 465211 48179 465277 48180
rect 465947 48244 466013 48245
rect 465947 48180 465948 48244
rect 466012 48180 466013 48244
rect 465947 48179 466013 48180
rect 466315 48244 466381 48245
rect 466315 48180 466316 48244
rect 466380 48180 466381 48244
rect 466315 48179 466381 48180
rect 467603 48244 467669 48245
rect 467603 48180 467604 48244
rect 467668 48180 467669 48244
rect 467603 48179 467669 48180
rect 468339 48244 468405 48245
rect 468339 48180 468340 48244
rect 468404 48180 468405 48244
rect 468339 48179 468405 48180
rect 468707 48244 468773 48245
rect 468707 48180 468708 48244
rect 468772 48180 468773 48244
rect 468707 48179 468773 48180
rect 469811 48244 469877 48245
rect 469811 48180 469812 48244
rect 469876 48180 469877 48244
rect 469811 48179 469877 48180
rect 470915 48244 470981 48245
rect 470915 48180 470916 48244
rect 470980 48180 470981 48244
rect 470915 48179 470981 48180
rect 471283 48244 471349 48245
rect 471283 48180 471284 48244
rect 471348 48180 471349 48244
rect 471283 48179 471349 48180
rect 472203 48244 472269 48245
rect 472203 48180 472204 48244
rect 472268 48180 472269 48244
rect 472203 48179 472269 48180
rect 460611 47700 460677 47701
rect 460611 47636 460612 47700
rect 460676 47636 460677 47700
rect 460611 47635 460677 47636
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 39454 470414 47940
rect 473310 47837 473370 49270
rect 474414 48245 474474 49950
rect 475702 49950 475828 50010
rect 475702 48245 475762 49950
rect 476040 49330 476100 50106
rect 476992 50010 477052 50106
rect 475886 49270 476100 49330
rect 476990 49950 477052 50010
rect 478080 50010 478140 50106
rect 478080 49950 478154 50010
rect 474411 48244 474477 48245
rect 474411 48180 474412 48244
rect 474476 48180 474477 48244
rect 474411 48179 474477 48180
rect 475699 48244 475765 48245
rect 475699 48180 475700 48244
rect 475764 48180 475765 48244
rect 475699 48179 475765 48180
rect 475886 47973 475946 49270
rect 476990 48245 477050 49950
rect 478094 48245 478154 49950
rect 478488 49877 478548 50106
rect 479168 50010 479228 50106
rect 479168 49950 479258 50010
rect 478485 49876 478551 49877
rect 478485 49812 478486 49876
rect 478550 49812 478551 49876
rect 478485 49811 478551 49812
rect 476987 48244 477053 48245
rect 476987 48180 476988 48244
rect 477052 48180 477053 48244
rect 476987 48179 477053 48180
rect 478091 48244 478157 48245
rect 478091 48180 478092 48244
rect 478156 48180 478157 48244
rect 478091 48179 478157 48180
rect 475883 47972 475949 47973
rect 473307 47836 473373 47837
rect 473307 47772 473308 47836
rect 473372 47772 473373 47836
rect 473307 47771 473373 47772
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 43174 474134 47940
rect 475883 47908 475884 47972
rect 475948 47908 475949 47972
rect 475883 47907 475949 47908
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 46894 477854 48064
rect 479198 47701 479258 49950
rect 480936 49877 480996 50106
rect 483520 50010 483580 50106
rect 483430 49950 483580 50010
rect 485968 50010 486028 50106
rect 485968 49950 486066 50010
rect 480933 49876 480999 49877
rect 480933 49812 480934 49876
rect 480998 49812 480999 49876
rect 480933 49811 480999 49812
rect 483430 49333 483490 49950
rect 486006 49469 486066 49950
rect 488280 49741 488340 50106
rect 488277 49740 488343 49741
rect 488277 49676 488278 49740
rect 488342 49676 488343 49740
rect 488277 49675 488343 49676
rect 491000 49605 491060 50106
rect 493448 49605 493508 50106
rect 495896 49741 495956 50106
rect 495893 49740 495959 49741
rect 495893 49676 495894 49740
rect 495958 49676 495959 49740
rect 495893 49675 495959 49676
rect 498480 49605 498540 50106
rect 500928 49605 500988 50106
rect 503512 49741 503572 50106
rect 503509 49740 503575 49741
rect 503509 49676 503510 49740
rect 503574 49676 503575 49740
rect 503509 49675 503575 49676
rect 505960 49605 506020 50106
rect 508544 49605 508604 50106
rect 510992 49605 511052 50106
rect 513440 49605 513500 50106
rect 515888 49605 515948 50106
rect 518472 50010 518532 50106
rect 518390 49950 518532 50010
rect 490997 49604 491063 49605
rect 490997 49540 490998 49604
rect 491062 49540 491063 49604
rect 490997 49539 491063 49540
rect 493445 49604 493511 49605
rect 493445 49540 493446 49604
rect 493510 49540 493511 49604
rect 493445 49539 493511 49540
rect 498477 49604 498543 49605
rect 498477 49540 498478 49604
rect 498542 49540 498543 49604
rect 498477 49539 498543 49540
rect 500925 49604 500991 49605
rect 500925 49540 500926 49604
rect 500990 49540 500991 49604
rect 500925 49539 500991 49540
rect 505957 49604 506023 49605
rect 505957 49540 505958 49604
rect 506022 49540 506023 49604
rect 505957 49539 506023 49540
rect 508541 49604 508607 49605
rect 508541 49540 508542 49604
rect 508606 49540 508607 49604
rect 508541 49539 508607 49540
rect 510989 49604 511055 49605
rect 510989 49540 510990 49604
rect 511054 49540 511055 49604
rect 510989 49539 511055 49540
rect 513437 49604 513503 49605
rect 513437 49540 513438 49604
rect 513502 49540 513503 49604
rect 513437 49539 513503 49540
rect 515885 49604 515951 49605
rect 515885 49540 515886 49604
rect 515950 49540 515951 49604
rect 515885 49539 515951 49540
rect 486003 49468 486069 49469
rect 486003 49404 486004 49468
rect 486068 49404 486069 49468
rect 486003 49403 486069 49404
rect 483427 49332 483493 49333
rect 483427 49268 483428 49332
rect 483492 49268 483493 49332
rect 483427 49267 483493 49268
rect 479195 47700 479261 47701
rect 479195 47636 479196 47700
rect 479260 47636 479261 47700
rect 479195 47635 479261 47636
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 14614 481574 47940
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 18334 485294 48064
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 22054 489014 47940
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 25774 492734 48064
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 29494 496454 47940
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 39454 506414 47940
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 43174 510134 48064
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 46894 513854 47940
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 14614 517574 48064
rect 518390 47157 518450 49950
rect 520920 49605 520980 50106
rect 523368 50010 523428 50106
rect 523358 49950 523428 50010
rect 520917 49604 520983 49605
rect 520917 49540 520918 49604
rect 520982 49540 520983 49604
rect 520917 49539 520983 49540
rect 518387 47156 518453 47157
rect 518387 47092 518388 47156
rect 518452 47092 518453 47156
rect 518387 47091 518453 47092
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 18334 521294 47940
rect 523358 47293 523418 49950
rect 525952 49605 526012 50106
rect 525949 49604 526015 49605
rect 525949 49540 525950 49604
rect 526014 49540 526015 49604
rect 525949 49539 526015 49540
rect 523355 47292 523421 47293
rect 523355 47228 523356 47292
rect 523420 47228 523421 47292
rect 523355 47227 523421 47228
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 22054 525014 48064
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 25774 528734 48064
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 29494 532454 48064
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 39454 542414 48064
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 43174 546134 48064
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 46894 549854 48064
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 48064
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 48064
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 60146 601538 60382 601774
rect 60466 601538 60702 601774
rect 60146 601218 60382 601454
rect 60466 601218 60702 601454
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 60146 565538 60382 565774
rect 60466 565538 60702 565774
rect 60146 565218 60382 565454
rect 60466 565218 60702 565454
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 63866 497258 64102 497494
rect 64186 497258 64422 497494
rect 63866 496938 64102 497174
rect 64186 496938 64422 497174
rect 63866 461258 64102 461494
rect 64186 461258 64422 461494
rect 63866 460938 64102 461174
rect 64186 460938 64422 461174
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 88706 486098 88942 486334
rect 89026 486098 89262 486334
rect 88706 485778 88942 486014
rect 89026 485778 89262 486014
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 92426 489818 92662 490054
rect 92746 489818 92982 490054
rect 92426 489498 92662 489734
rect 92746 489498 92982 489734
rect 92426 453818 92662 454054
rect 92746 453818 92982 454054
rect 92426 453498 92662 453734
rect 92746 453498 92982 453734
rect 96146 493538 96382 493774
rect 96466 493538 96702 493774
rect 96146 493218 96382 493454
rect 96466 493218 96702 493454
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 99866 497258 100102 497494
rect 100186 497258 100422 497494
rect 99866 496938 100102 497174
rect 100186 496938 100422 497174
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 128426 489818 128662 490054
rect 128746 489818 128982 490054
rect 128426 489498 128662 489734
rect 128746 489498 128982 489734
rect 128426 453818 128662 454054
rect 128746 453818 128982 454054
rect 128426 453498 128662 453734
rect 128746 453498 128982 453734
rect 132146 493538 132382 493774
rect 132466 493538 132702 493774
rect 132146 493218 132382 493454
rect 132466 493218 132702 493454
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 135866 497258 136102 497494
rect 136186 497258 136422 497494
rect 135866 496938 136102 497174
rect 136186 496938 136422 497174
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 164426 597818 164662 598054
rect 164746 597818 164982 598054
rect 164426 597498 164662 597734
rect 164746 597498 164982 597734
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 164426 561818 164662 562054
rect 164746 561818 164982 562054
rect 164426 561498 164662 561734
rect 164746 561498 164982 561734
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 164426 525818 164662 526054
rect 164746 525818 164982 526054
rect 164426 525498 164662 525734
rect 164746 525498 164982 525734
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 160706 486098 160942 486334
rect 161026 486098 161262 486334
rect 160706 485778 160942 486014
rect 161026 485778 161262 486014
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 160706 414098 160942 414334
rect 161026 414098 161262 414334
rect 160706 413778 160942 414014
rect 161026 413778 161262 414014
rect 20328 402938 20564 403174
rect 20328 402618 20564 402854
rect 156056 402938 156292 403174
rect 156056 402618 156292 402854
rect 21008 399218 21244 399454
rect 21008 398898 21244 399134
rect 155376 399218 155612 399454
rect 155376 398898 155612 399134
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 20328 366938 20564 367174
rect 20328 366618 20564 366854
rect 156056 366938 156292 367174
rect 156056 366618 156292 366854
rect 21008 363218 21244 363454
rect 21008 362898 21244 363134
rect 155376 363218 155612 363454
rect 155376 362898 155612 363134
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 20328 330938 20564 331174
rect 20328 330618 20564 330854
rect 156056 330938 156292 331174
rect 156056 330618 156292 330854
rect 21008 327218 21244 327454
rect 21008 326898 21244 327134
rect 155376 327218 155612 327454
rect 155376 326898 155612 327134
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 20328 294938 20564 295174
rect 20328 294618 20564 294854
rect 156056 294938 156292 295174
rect 156056 294618 156292 294854
rect 21008 291218 21244 291454
rect 21008 290898 21244 291134
rect 155376 291218 155612 291454
rect 155376 290898 155612 291134
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 20328 258938 20564 259174
rect 20328 258618 20564 258854
rect 156056 258938 156292 259174
rect 156056 258618 156292 258854
rect 21008 255218 21244 255454
rect 21008 254898 21244 255134
rect 155376 255218 155612 255454
rect 155376 254898 155612 255134
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 20328 222938 20564 223174
rect 20328 222618 20564 222854
rect 156056 222938 156292 223174
rect 156056 222618 156292 222854
rect 21008 219218 21244 219454
rect 21008 218898 21244 219134
rect 155376 219218 155612 219454
rect 155376 218898 155612 219134
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 20328 186938 20564 187174
rect 20328 186618 20564 186854
rect 156056 186938 156292 187174
rect 156056 186618 156292 186854
rect 21008 183218 21244 183454
rect 21008 182898 21244 183134
rect 155376 183218 155612 183454
rect 155376 182898 155612 183134
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 20328 150938 20564 151174
rect 20328 150618 20564 150854
rect 156056 150938 156292 151174
rect 156056 150618 156292 150854
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 20328 114938 20564 115174
rect 20328 114618 20564 114854
rect 156056 114938 156292 115174
rect 156056 114618 156292 114854
rect 21008 111218 21244 111454
rect 21008 110898 21244 111134
rect 155376 111218 155612 111454
rect 155376 110898 155612 111134
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 20328 78938 20564 79174
rect 20328 78618 20564 78854
rect 156056 78938 156292 79174
rect 156056 78618 156292 78854
rect 21008 75218 21244 75454
rect 21008 74898 21244 75134
rect 155376 75218 155612 75454
rect 155376 74898 155612 75134
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 489818 164662 490054
rect 164746 489818 164982 490054
rect 164426 489498 164662 489734
rect 164746 489498 164982 489734
rect 164426 453818 164662 454054
rect 164746 453818 164982 454054
rect 164426 453498 164662 453734
rect 164746 453498 164982 453734
rect 164426 417818 164662 418054
rect 164746 417818 164982 418054
rect 164426 417498 164662 417734
rect 164746 417498 164982 417734
rect 164426 381818 164662 382054
rect 164746 381818 164982 382054
rect 164426 381498 164662 381734
rect 164746 381498 164982 381734
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 168146 493538 168382 493774
rect 168466 493538 168702 493774
rect 168146 493218 168382 493454
rect 168466 493218 168702 493454
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 168146 421538 168382 421774
rect 168466 421538 168702 421774
rect 168146 421218 168382 421454
rect 168466 421218 168702 421454
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 171866 497258 172102 497494
rect 172186 497258 172422 497494
rect 171866 496938 172102 497174
rect 172186 496938 172422 497174
rect 171866 461258 172102 461494
rect 172186 461258 172422 461494
rect 171866 460938 172102 461174
rect 172186 460938 172422 461174
rect 171866 425258 172102 425494
rect 172186 425258 172422 425494
rect 171866 424938 172102 425174
rect 172186 424938 172422 425174
rect 171866 389258 172102 389494
rect 172186 389258 172422 389494
rect 171866 388938 172102 389174
rect 172186 388938 172422 389174
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 196706 594098 196942 594334
rect 197026 594098 197262 594334
rect 196706 593778 196942 594014
rect 197026 593778 197262 594014
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 194250 435218 194486 435454
rect 194250 434898 194486 435134
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 194250 399218 194486 399454
rect 194250 398898 194486 399134
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 194250 363218 194486 363454
rect 194250 362898 194486 363134
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 194250 327218 194486 327454
rect 194250 326898 194486 327134
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 194250 291218 194486 291454
rect 194250 290898 194486 291134
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 194250 255218 194486 255454
rect 194250 254898 194486 255134
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 200426 597818 200662 598054
rect 200746 597818 200982 598054
rect 200426 597498 200662 597734
rect 200746 597498 200982 597734
rect 200426 561818 200662 562054
rect 200746 561818 200982 562054
rect 200426 561498 200662 561734
rect 200746 561498 200982 561734
rect 200426 525818 200662 526054
rect 200746 525818 200982 526054
rect 200426 525498 200662 525734
rect 200746 525498 200982 525734
rect 200426 489818 200662 490054
rect 200746 489818 200982 490054
rect 200426 489498 200662 489734
rect 200746 489498 200982 489734
rect 200426 453818 200662 454054
rect 200746 453818 200982 454054
rect 200426 453498 200662 453734
rect 200746 453498 200982 453734
rect 200426 417818 200662 418054
rect 200746 417818 200982 418054
rect 200426 417498 200662 417734
rect 200746 417498 200982 417734
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 200426 273818 200662 274054
rect 200746 273818 200982 274054
rect 200426 273498 200662 273734
rect 200746 273498 200982 273734
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 200426 201818 200662 202054
rect 200746 201818 200982 202054
rect 200426 201498 200662 201734
rect 200746 201498 200982 201734
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 204146 601538 204382 601774
rect 204466 601538 204702 601774
rect 204146 601218 204382 601454
rect 204466 601218 204702 601454
rect 204146 565538 204382 565774
rect 204466 565538 204702 565774
rect 204146 565218 204382 565454
rect 204466 565218 204702 565454
rect 204146 529538 204382 529774
rect 204466 529538 204702 529774
rect 204146 529218 204382 529454
rect 204466 529218 204702 529454
rect 204146 493538 204382 493774
rect 204466 493538 204702 493774
rect 204146 493218 204382 493454
rect 204466 493218 204702 493454
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 204146 421538 204382 421774
rect 204466 421538 204702 421774
rect 204146 421218 204382 421454
rect 204466 421218 204702 421454
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 207866 605258 208102 605494
rect 208186 605258 208422 605494
rect 207866 604938 208102 605174
rect 208186 604938 208422 605174
rect 207866 569258 208102 569494
rect 208186 569258 208422 569494
rect 207866 568938 208102 569174
rect 208186 568938 208422 569174
rect 207866 533258 208102 533494
rect 208186 533258 208422 533494
rect 207866 532938 208102 533174
rect 208186 532938 208422 533174
rect 207866 497258 208102 497494
rect 208186 497258 208422 497494
rect 207866 496938 208102 497174
rect 208186 496938 208422 497174
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 209610 438938 209846 439174
rect 209610 438618 209846 438854
rect 207866 425258 208102 425494
rect 208186 425258 208422 425494
rect 207866 424938 208102 425174
rect 208186 424938 208422 425174
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 209610 402938 209846 403174
rect 209610 402618 209846 402854
rect 207866 389258 208102 389494
rect 208186 389258 208422 389494
rect 207866 388938 208102 389174
rect 208186 388938 208422 389174
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 209610 366938 209846 367174
rect 209610 366618 209846 366854
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 209610 330938 209846 331174
rect 209610 330618 209846 330854
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 209610 294938 209846 295174
rect 209610 294618 209846 294854
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 209610 258938 209846 259174
rect 209610 258618 209846 258854
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 224970 435218 225206 435454
rect 224970 434898 225206 435134
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 224970 399218 225206 399454
rect 224970 398898 225206 399134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 224970 363218 225206 363454
rect 224970 362898 225206 363134
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 224970 327218 225206 327454
rect 224970 326898 225206 327134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 224970 291218 225206 291454
rect 224970 290898 225206 291134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 224970 255218 225206 255454
rect 224970 254898 225206 255134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 232706 630098 232942 630334
rect 233026 630098 233262 630334
rect 232706 629778 232942 630014
rect 233026 629778 233262 630014
rect 232706 594098 232942 594334
rect 233026 594098 233262 594334
rect 232706 593778 232942 594014
rect 233026 593778 233262 594014
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 232706 522098 232942 522334
rect 233026 522098 233262 522334
rect 232706 521778 232942 522014
rect 233026 521778 233262 522014
rect 232706 486098 232942 486334
rect 233026 486098 233262 486334
rect 232706 485778 232942 486014
rect 233026 485778 233262 486014
rect 232706 450098 232942 450334
rect 233026 450098 233262 450334
rect 232706 449778 232942 450014
rect 233026 449778 233262 450014
rect 232706 414098 232942 414334
rect 233026 414098 233262 414334
rect 232706 413778 232942 414014
rect 233026 413778 233262 414014
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 236426 597818 236662 598054
rect 236746 597818 236982 598054
rect 236426 597498 236662 597734
rect 236746 597498 236982 597734
rect 236426 561818 236662 562054
rect 236746 561818 236982 562054
rect 236426 561498 236662 561734
rect 236746 561498 236982 561734
rect 236426 525818 236662 526054
rect 236746 525818 236982 526054
rect 236426 525498 236662 525734
rect 236746 525498 236982 525734
rect 236426 489818 236662 490054
rect 236746 489818 236982 490054
rect 236426 489498 236662 489734
rect 236746 489498 236982 489734
rect 236426 453818 236662 454054
rect 236746 453818 236982 454054
rect 236426 453498 236662 453734
rect 236746 453498 236982 453734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 240146 601538 240382 601774
rect 240466 601538 240702 601774
rect 240146 601218 240382 601454
rect 240466 601218 240702 601454
rect 240146 565538 240382 565774
rect 240466 565538 240702 565774
rect 240146 565218 240382 565454
rect 240466 565218 240702 565454
rect 240146 529538 240382 529774
rect 240466 529538 240702 529774
rect 240146 529218 240382 529454
rect 240466 529218 240702 529454
rect 240146 493538 240382 493774
rect 240466 493538 240702 493774
rect 240146 493218 240382 493454
rect 240466 493218 240702 493454
rect 240146 457538 240382 457774
rect 240466 457538 240702 457774
rect 240146 457218 240382 457454
rect 240466 457218 240702 457454
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 243866 605258 244102 605494
rect 244186 605258 244422 605494
rect 243866 604938 244102 605174
rect 244186 604938 244422 605174
rect 243866 569258 244102 569494
rect 244186 569258 244422 569494
rect 243866 568938 244102 569174
rect 244186 568938 244422 569174
rect 243866 533258 244102 533494
rect 244186 533258 244422 533494
rect 243866 532938 244102 533174
rect 244186 532938 244422 533174
rect 243866 497258 244102 497494
rect 244186 497258 244422 497494
rect 243866 496938 244102 497174
rect 244186 496938 244422 497174
rect 243866 461258 244102 461494
rect 244186 461258 244422 461494
rect 243866 460938 244102 461174
rect 244186 460938 244422 461174
rect 240330 438938 240566 439174
rect 240330 438618 240566 438854
rect 236426 417818 236662 418054
rect 236746 417818 236982 418054
rect 236426 417498 236662 417734
rect 236746 417498 236982 417734
rect 243866 425258 244102 425494
rect 244186 425258 244422 425494
rect 243866 424938 244102 425174
rect 244186 424938 244422 425174
rect 240330 402938 240566 403174
rect 240330 402618 240566 402854
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 243866 389258 244102 389494
rect 244186 389258 244422 389494
rect 243866 388938 244102 389174
rect 244186 388938 244422 389174
rect 240330 366938 240566 367174
rect 240330 366618 240566 366854
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 243866 353258 244102 353494
rect 244186 353258 244422 353494
rect 243866 352938 244102 353174
rect 244186 352938 244422 353174
rect 240330 330938 240566 331174
rect 240330 330618 240566 330854
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 243866 317258 244102 317494
rect 244186 317258 244422 317494
rect 243866 316938 244102 317174
rect 244186 316938 244422 317174
rect 240330 294938 240566 295174
rect 240330 294618 240566 294854
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 243866 281258 244102 281494
rect 244186 281258 244422 281494
rect 243866 280938 244102 281174
rect 244186 280938 244422 281174
rect 240330 258938 240566 259174
rect 240330 258618 240566 258854
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 236426 93818 236662 94054
rect 236746 93818 236982 94054
rect 236426 93498 236662 93734
rect 236746 93498 236982 93734
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 241538 240382 241774
rect 240466 241538 240702 241774
rect 240146 241218 240382 241454
rect 240466 241218 240702 241454
rect 240146 205538 240382 205774
rect 240466 205538 240702 205774
rect 240146 205218 240382 205454
rect 240466 205218 240702 205454
rect 240146 169538 240382 169774
rect 240466 169538 240702 169774
rect 240146 169218 240382 169454
rect 240466 169218 240702 169454
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 245258 244102 245494
rect 244186 245258 244422 245494
rect 243866 244938 244102 245174
rect 244186 244938 244422 245174
rect 243866 209258 244102 209494
rect 244186 209258 244422 209494
rect 243866 208938 244102 209174
rect 244186 208938 244422 209174
rect 243866 173258 244102 173494
rect 244186 173258 244422 173494
rect 243866 172938 244102 173174
rect 244186 172938 244422 173174
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 268706 630098 268942 630334
rect 269026 630098 269262 630334
rect 268706 629778 268942 630014
rect 269026 629778 269262 630014
rect 268706 594098 268942 594334
rect 269026 594098 269262 594334
rect 268706 593778 268942 594014
rect 269026 593778 269262 594014
rect 268706 558098 268942 558334
rect 269026 558098 269262 558334
rect 268706 557778 268942 558014
rect 269026 557778 269262 558014
rect 268706 522098 268942 522334
rect 269026 522098 269262 522334
rect 268706 521778 268942 522014
rect 269026 521778 269262 522014
rect 268706 486098 268942 486334
rect 269026 486098 269262 486334
rect 268706 485778 268942 486014
rect 269026 485778 269262 486014
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 272426 633818 272662 634054
rect 272746 633818 272982 634054
rect 272426 633498 272662 633734
rect 272746 633498 272982 633734
rect 272426 597818 272662 598054
rect 272746 597818 272982 598054
rect 272426 597498 272662 597734
rect 272746 597498 272982 597734
rect 272426 561818 272662 562054
rect 272746 561818 272982 562054
rect 272426 561498 272662 561734
rect 272746 561498 272982 561734
rect 272426 525818 272662 526054
rect 272746 525818 272982 526054
rect 272426 525498 272662 525734
rect 272746 525498 272982 525734
rect 272426 489818 272662 490054
rect 272746 489818 272982 490054
rect 272426 489498 272662 489734
rect 272746 489498 272982 489734
rect 272426 453818 272662 454054
rect 272746 453818 272982 454054
rect 272426 453498 272662 453734
rect 272746 453498 272982 453734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 276146 637538 276382 637774
rect 276466 637538 276702 637774
rect 276146 637218 276382 637454
rect 276466 637218 276702 637454
rect 276146 601538 276382 601774
rect 276466 601538 276702 601774
rect 276146 601218 276382 601454
rect 276466 601218 276702 601454
rect 276146 565538 276382 565774
rect 276466 565538 276702 565774
rect 276146 565218 276382 565454
rect 276466 565218 276702 565454
rect 276146 529538 276382 529774
rect 276466 529538 276702 529774
rect 276146 529218 276382 529454
rect 276466 529218 276702 529454
rect 276146 493538 276382 493774
rect 276466 493538 276702 493774
rect 276146 493218 276382 493454
rect 276466 493218 276702 493454
rect 276146 457538 276382 457774
rect 276466 457538 276702 457774
rect 276146 457218 276382 457454
rect 276466 457218 276702 457454
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 279866 641258 280102 641494
rect 280186 641258 280422 641494
rect 279866 640938 280102 641174
rect 280186 640938 280422 641174
rect 279866 605258 280102 605494
rect 280186 605258 280422 605494
rect 279866 604938 280102 605174
rect 280186 604938 280422 605174
rect 279866 569258 280102 569494
rect 280186 569258 280422 569494
rect 279866 568938 280102 569174
rect 280186 568938 280422 569174
rect 279866 533258 280102 533494
rect 280186 533258 280422 533494
rect 279866 532938 280102 533174
rect 280186 532938 280422 533174
rect 279866 497258 280102 497494
rect 280186 497258 280422 497494
rect 279866 496938 280102 497174
rect 280186 496938 280422 497174
rect 279866 461258 280102 461494
rect 280186 461258 280422 461494
rect 279866 460938 280102 461174
rect 280186 460938 280422 461174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 304706 630098 304942 630334
rect 305026 630098 305262 630334
rect 304706 629778 304942 630014
rect 305026 629778 305262 630014
rect 304706 594098 304942 594334
rect 305026 594098 305262 594334
rect 304706 593778 304942 594014
rect 305026 593778 305262 594014
rect 304706 558098 304942 558334
rect 305026 558098 305262 558334
rect 304706 557778 304942 558014
rect 305026 557778 305262 558014
rect 304706 522098 304942 522334
rect 305026 522098 305262 522334
rect 304706 521778 304942 522014
rect 305026 521778 305262 522014
rect 304706 486098 304942 486334
rect 305026 486098 305262 486334
rect 304706 485778 304942 486014
rect 305026 485778 305262 486014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 308426 633818 308662 634054
rect 308746 633818 308982 634054
rect 308426 633498 308662 633734
rect 308746 633498 308982 633734
rect 308426 597818 308662 598054
rect 308746 597818 308982 598054
rect 308426 597498 308662 597734
rect 308746 597498 308982 597734
rect 308426 561818 308662 562054
rect 308746 561818 308982 562054
rect 308426 561498 308662 561734
rect 308746 561498 308982 561734
rect 308426 525818 308662 526054
rect 308746 525818 308982 526054
rect 308426 525498 308662 525734
rect 308746 525498 308982 525734
rect 308426 489818 308662 490054
rect 308746 489818 308982 490054
rect 308426 489498 308662 489734
rect 308746 489498 308982 489734
rect 308426 453818 308662 454054
rect 308746 453818 308982 454054
rect 308426 453498 308662 453734
rect 308746 453498 308982 453734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 312146 637538 312382 637774
rect 312466 637538 312702 637774
rect 312146 637218 312382 637454
rect 312466 637218 312702 637454
rect 312146 601538 312382 601774
rect 312466 601538 312702 601774
rect 312146 601218 312382 601454
rect 312466 601218 312702 601454
rect 312146 565538 312382 565774
rect 312466 565538 312702 565774
rect 312146 565218 312382 565454
rect 312466 565218 312702 565454
rect 312146 529538 312382 529774
rect 312466 529538 312702 529774
rect 312146 529218 312382 529454
rect 312466 529218 312702 529454
rect 312146 493538 312382 493774
rect 312466 493538 312702 493774
rect 312146 493218 312382 493454
rect 312466 493218 312702 493454
rect 312146 457538 312382 457774
rect 312466 457538 312702 457774
rect 312146 457218 312382 457454
rect 312466 457218 312702 457454
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 315866 641258 316102 641494
rect 316186 641258 316422 641494
rect 315866 640938 316102 641174
rect 316186 640938 316422 641174
rect 315866 605258 316102 605494
rect 316186 605258 316422 605494
rect 315866 604938 316102 605174
rect 316186 604938 316422 605174
rect 315866 569258 316102 569494
rect 316186 569258 316422 569494
rect 315866 568938 316102 569174
rect 316186 568938 316422 569174
rect 315866 533258 316102 533494
rect 316186 533258 316422 533494
rect 315866 532938 316102 533174
rect 316186 532938 316422 533174
rect 315866 497258 316102 497494
rect 316186 497258 316422 497494
rect 315866 496938 316102 497174
rect 316186 496938 316422 497174
rect 315866 461258 316102 461494
rect 316186 461258 316422 461494
rect 315866 460938 316102 461174
rect 316186 460938 316422 461174
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 340706 630098 340942 630334
rect 341026 630098 341262 630334
rect 340706 629778 340942 630014
rect 341026 629778 341262 630014
rect 340706 594098 340942 594334
rect 341026 594098 341262 594334
rect 340706 593778 340942 594014
rect 341026 593778 341262 594014
rect 340706 558098 340942 558334
rect 341026 558098 341262 558334
rect 340706 557778 340942 558014
rect 341026 557778 341262 558014
rect 340706 522098 340942 522334
rect 341026 522098 341262 522334
rect 340706 521778 340942 522014
rect 341026 521778 341262 522014
rect 340706 486098 340942 486334
rect 341026 486098 341262 486334
rect 340706 485778 340942 486014
rect 341026 485778 341262 486014
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 344426 597818 344662 598054
rect 344746 597818 344982 598054
rect 344426 597498 344662 597734
rect 344746 597498 344982 597734
rect 344426 561818 344662 562054
rect 344746 561818 344982 562054
rect 344426 561498 344662 561734
rect 344746 561498 344982 561734
rect 344426 525818 344662 526054
rect 344746 525818 344982 526054
rect 344426 525498 344662 525734
rect 344746 525498 344982 525734
rect 344426 489818 344662 490054
rect 344746 489818 344982 490054
rect 344426 489498 344662 489734
rect 344746 489498 344982 489734
rect 344426 453818 344662 454054
rect 344746 453818 344982 454054
rect 344426 453498 344662 453734
rect 344746 453498 344982 453734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 348146 601538 348382 601774
rect 348466 601538 348702 601774
rect 348146 601218 348382 601454
rect 348466 601218 348702 601454
rect 348146 565538 348382 565774
rect 348466 565538 348702 565774
rect 348146 565218 348382 565454
rect 348466 565218 348702 565454
rect 348146 529538 348382 529774
rect 348466 529538 348702 529774
rect 348146 529218 348382 529454
rect 348466 529218 348702 529454
rect 348146 493538 348382 493774
rect 348466 493538 348702 493774
rect 348146 493218 348382 493454
rect 348466 493218 348702 493454
rect 348146 457538 348382 457774
rect 348466 457538 348702 457774
rect 348146 457218 348382 457454
rect 348466 457218 348702 457454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 351866 605258 352102 605494
rect 352186 605258 352422 605494
rect 351866 604938 352102 605174
rect 352186 604938 352422 605174
rect 351866 569258 352102 569494
rect 352186 569258 352422 569494
rect 351866 568938 352102 569174
rect 352186 568938 352422 569174
rect 351866 533258 352102 533494
rect 352186 533258 352422 533494
rect 351866 532938 352102 533174
rect 352186 532938 352422 533174
rect 351866 497258 352102 497494
rect 352186 497258 352422 497494
rect 351866 496938 352102 497174
rect 352186 496938 352422 497174
rect 351866 461258 352102 461494
rect 352186 461258 352422 461494
rect 351866 460938 352102 461174
rect 352186 460938 352422 461174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 271050 438938 271286 439174
rect 271050 438618 271286 438854
rect 301770 438938 302006 439174
rect 301770 438618 302006 438854
rect 332490 438938 332726 439174
rect 332490 438618 332726 438854
rect 363210 438938 363446 439174
rect 363210 438618 363446 438854
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 255690 435218 255926 435454
rect 255690 434898 255926 435134
rect 286410 435218 286646 435454
rect 286410 434898 286646 435134
rect 317130 435218 317366 435454
rect 317130 434898 317366 435134
rect 347850 435218 348086 435454
rect 347850 434898 348086 435134
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 271050 402938 271286 403174
rect 271050 402618 271286 402854
rect 301770 402938 302006 403174
rect 301770 402618 302006 402854
rect 332490 402938 332726 403174
rect 332490 402618 332726 402854
rect 363210 402938 363446 403174
rect 363210 402618 363446 402854
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 255690 399218 255926 399454
rect 255690 398898 255926 399134
rect 286410 399218 286646 399454
rect 286410 398898 286646 399134
rect 317130 399218 317366 399454
rect 317130 398898 317366 399134
rect 347850 399218 348086 399454
rect 347850 398898 348086 399134
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 271050 366938 271286 367174
rect 271050 366618 271286 366854
rect 301770 366938 302006 367174
rect 301770 366618 302006 366854
rect 332490 366938 332726 367174
rect 332490 366618 332726 366854
rect 363210 366938 363446 367174
rect 363210 366618 363446 366854
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 255690 363218 255926 363454
rect 255690 362898 255926 363134
rect 286410 363218 286646 363454
rect 286410 362898 286646 363134
rect 317130 363218 317366 363454
rect 317130 362898 317366 363134
rect 347850 363218 348086 363454
rect 347850 362898 348086 363134
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 271050 330938 271286 331174
rect 271050 330618 271286 330854
rect 301770 330938 302006 331174
rect 301770 330618 302006 330854
rect 332490 330938 332726 331174
rect 332490 330618 332726 330854
rect 363210 330938 363446 331174
rect 363210 330618 363446 330854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 255690 327218 255926 327454
rect 255690 326898 255926 327134
rect 286410 327218 286646 327454
rect 286410 326898 286646 327134
rect 317130 327218 317366 327454
rect 317130 326898 317366 327134
rect 347850 327218 348086 327454
rect 347850 326898 348086 327134
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 271050 294938 271286 295174
rect 271050 294618 271286 294854
rect 301770 294938 302006 295174
rect 301770 294618 302006 294854
rect 332490 294938 332726 295174
rect 332490 294618 332726 294854
rect 363210 294938 363446 295174
rect 363210 294618 363446 294854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 255690 291218 255926 291454
rect 255690 290898 255926 291134
rect 286410 291218 286646 291454
rect 286410 290898 286646 291134
rect 317130 291218 317366 291454
rect 317130 290898 317366 291134
rect 347850 291218 348086 291454
rect 347850 290898 348086 291134
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 271050 258938 271286 259174
rect 271050 258618 271286 258854
rect 301770 258938 302006 259174
rect 301770 258618 302006 258854
rect 332490 258938 332726 259174
rect 332490 258618 332726 258854
rect 363210 258938 363446 259174
rect 363210 258618 363446 258854
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 255690 255218 255926 255454
rect 255690 254898 255926 255134
rect 286410 255218 286646 255454
rect 286410 254898 286646 255134
rect 317130 255218 317366 255454
rect 317130 254898 317366 255134
rect 347850 255218 348086 255454
rect 347850 254898 348086 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 234098 268942 234334
rect 269026 234098 269262 234334
rect 268706 233778 268942 234014
rect 269026 233778 269262 234014
rect 268706 198098 268942 198334
rect 269026 198098 269262 198334
rect 268706 197778 268942 198014
rect 269026 197778 269262 198014
rect 268706 162098 268942 162334
rect 269026 162098 269262 162334
rect 268706 161778 268942 162014
rect 269026 161778 269262 162014
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 268706 90098 268942 90334
rect 269026 90098 269262 90334
rect 268706 89778 268942 90014
rect 269026 89778 269262 90014
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 237818 272662 238054
rect 272746 237818 272982 238054
rect 272426 237498 272662 237734
rect 272746 237498 272982 237734
rect 272426 201818 272662 202054
rect 272746 201818 272982 202054
rect 272426 201498 272662 201734
rect 272746 201498 272982 201734
rect 272426 165818 272662 166054
rect 272746 165818 272982 166054
rect 272426 165498 272662 165734
rect 272746 165498 272982 165734
rect 272426 129818 272662 130054
rect 272746 129818 272982 130054
rect 272426 129498 272662 129734
rect 272746 129498 272982 129734
rect 272426 93818 272662 94054
rect 272746 93818 272982 94054
rect 272426 93498 272662 93734
rect 272746 93498 272982 93734
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 241538 276382 241774
rect 276466 241538 276702 241774
rect 276146 241218 276382 241454
rect 276466 241218 276702 241454
rect 276146 205538 276382 205774
rect 276466 205538 276702 205774
rect 276146 205218 276382 205454
rect 276466 205218 276702 205454
rect 276146 169538 276382 169774
rect 276466 169538 276702 169774
rect 276146 169218 276382 169454
rect 276466 169218 276702 169454
rect 276146 133538 276382 133774
rect 276466 133538 276702 133774
rect 276146 133218 276382 133454
rect 276466 133218 276702 133454
rect 276146 97538 276382 97774
rect 276466 97538 276702 97774
rect 276146 97218 276382 97454
rect 276466 97218 276702 97454
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 245258 280102 245494
rect 280186 245258 280422 245494
rect 279866 244938 280102 245174
rect 280186 244938 280422 245174
rect 279866 209258 280102 209494
rect 280186 209258 280422 209494
rect 279866 208938 280102 209174
rect 280186 208938 280422 209174
rect 279866 173258 280102 173494
rect 280186 173258 280422 173494
rect 279866 172938 280102 173174
rect 280186 172938 280422 173174
rect 279866 137258 280102 137494
rect 280186 137258 280422 137494
rect 279866 136938 280102 137174
rect 280186 136938 280422 137174
rect 279866 101258 280102 101494
rect 280186 101258 280422 101494
rect 279866 100938 280102 101174
rect 280186 100938 280422 101174
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 237818 308662 238054
rect 308746 237818 308982 238054
rect 308426 237498 308662 237734
rect 308746 237498 308982 237734
rect 308426 201818 308662 202054
rect 308746 201818 308982 202054
rect 308426 201498 308662 201734
rect 308746 201498 308982 201734
rect 308426 165818 308662 166054
rect 308746 165818 308982 166054
rect 308426 165498 308662 165734
rect 308746 165498 308982 165734
rect 308426 129818 308662 130054
rect 308746 129818 308982 130054
rect 308426 129498 308662 129734
rect 308746 129498 308982 129734
rect 308426 93818 308662 94054
rect 308746 93818 308982 94054
rect 308426 93498 308662 93734
rect 308746 93498 308982 93734
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 340706 90098 340942 90334
rect 341026 90098 341262 90334
rect 340706 89778 340942 90014
rect 341026 89778 341262 90014
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 378570 435218 378806 435454
rect 378570 434898 378806 435134
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 378570 399218 378806 399454
rect 378570 398898 378806 399134
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 378570 363218 378806 363454
rect 378570 362898 378806 363134
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 378570 327218 378806 327454
rect 378570 326898 378806 327134
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 378570 291218 378806 291454
rect 378570 290898 378806 291134
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 378570 255218 378806 255454
rect 378570 254898 378806 255134
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 459866 641258 460102 641494
rect 460186 641258 460422 641494
rect 459866 640938 460102 641174
rect 460186 640938 460422 641174
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 484706 630098 484942 630334
rect 485026 630098 485262 630334
rect 484706 629778 484942 630014
rect 485026 629778 485262 630014
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 488426 633818 488662 634054
rect 488746 633818 488982 634054
rect 488426 633498 488662 633734
rect 488746 633498 488982 633734
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 492146 637538 492382 637774
rect 492466 637538 492702 637774
rect 492146 637218 492382 637454
rect 492466 637218 492702 637454
rect 492146 601538 492382 601774
rect 492466 601538 492702 601774
rect 492146 601218 492382 601454
rect 492466 601218 492702 601454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 495866 641258 496102 641494
rect 496186 641258 496422 641494
rect 495866 640938 496102 641174
rect 496186 640938 496422 641174
rect 495866 605258 496102 605494
rect 496186 605258 496422 605494
rect 495866 604938 496102 605174
rect 496186 604938 496422 605174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 420328 582693 420564 582929
rect 556056 582693 556292 582929
rect 421008 579218 421244 579454
rect 421008 578898 421244 579134
rect 555376 579218 555612 579454
rect 555376 578898 555612 579134
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 420328 546938 420564 547174
rect 420328 546618 420564 546854
rect 556056 546938 556292 547174
rect 556056 546618 556292 546854
rect 421008 543218 421244 543454
rect 421008 542898 421244 543134
rect 555376 543218 555612 543454
rect 555376 542898 555612 543134
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 420328 510938 420564 511174
rect 420328 510618 420564 510854
rect 556056 510938 556292 511174
rect 556056 510618 556292 510854
rect 421008 507218 421244 507454
rect 421008 506898 421244 507134
rect 555376 507218 555612 507454
rect 555376 506898 555612 507134
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 420328 402938 420564 403174
rect 420328 402618 420564 402854
rect 556056 402938 556292 403174
rect 556056 402618 556292 402854
rect 421008 399218 421244 399454
rect 421008 398898 421244 399134
rect 555376 399218 555612 399454
rect 555376 398898 555612 399134
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 420328 366938 420564 367174
rect 420328 366618 420564 366854
rect 556056 366938 556292 367174
rect 556056 366618 556292 366854
rect 421008 363218 421244 363454
rect 421008 362898 421244 363134
rect 555376 363218 555612 363454
rect 555376 362898 555612 363134
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 420328 330938 420564 331174
rect 420328 330618 420564 330854
rect 556056 330938 556292 331174
rect 556056 330618 556292 330854
rect 421008 327218 421244 327454
rect 421008 326898 421244 327134
rect 555376 327218 555612 327454
rect 555376 326898 555612 327134
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 420328 294938 420564 295174
rect 420328 294618 420564 294854
rect 556056 294938 556292 295174
rect 556056 294618 556292 294854
rect 421008 291218 421244 291454
rect 421008 290898 421244 291134
rect 555376 291218 555612 291454
rect 555376 290898 555612 291134
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 420328 258938 420564 259174
rect 420328 258618 420564 258854
rect 556056 258938 556292 259174
rect 556056 258618 556292 258854
rect 421008 255218 421244 255454
rect 421008 254898 421244 255134
rect 555376 255218 555612 255454
rect 555376 254898 555612 255134
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 420328 222938 420564 223174
rect 420328 222618 420564 222854
rect 556056 222938 556292 223174
rect 556056 222618 556292 222854
rect 421008 219218 421244 219454
rect 421008 218898 421244 219134
rect 555376 219218 555612 219454
rect 555376 218898 555612 219134
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 420328 186938 420564 187174
rect 420328 186618 420564 186854
rect 556056 186938 556292 187174
rect 556056 186618 556292 186854
rect 421008 183218 421244 183454
rect 421008 182898 421244 183134
rect 555376 183218 555612 183454
rect 555376 182898 555612 183134
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 420328 150938 420564 151174
rect 420328 150618 420564 150854
rect 556056 150938 556292 151174
rect 556056 150618 556292 150854
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 420328 114938 420564 115174
rect 420328 114618 420564 114854
rect 556056 114938 556292 115174
rect 556056 114618 556292 114854
rect 421008 111218 421244 111454
rect 421008 110898 421244 111134
rect 555376 111218 555612 111454
rect 555376 110898 555612 111134
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 420328 78938 420564 79174
rect 420328 78618 420564 78854
rect 556056 78938 556292 79174
rect 556056 78618 556292 78854
rect 421008 75218 421244 75454
rect 421008 74898 421244 75134
rect 555376 75218 555612 75454
rect 555376 74898 555612 75134
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 193210 655174
rect 193446 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 193210 654854
rect 193446 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 495866 641494
rect 496102 641258 496186 641494
rect 496422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 495866 641174
rect 496102 640938 496186 641174
rect 496422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 193210 619174
rect 193446 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 193210 618854
rect 193446 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 495866 605494
rect 496102 605258 496186 605494
rect 496422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 495866 605174
rect 496102 604938 496186 605174
rect 496422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 193210 583174
rect 193446 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582929 592650 582938
rect -8726 582854 420328 582929
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 193210 582854
rect 193446 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582693 420328 582854
rect 420564 582693 556056 582929
rect 556292 582854 592650 582929
rect 556292 582693 581546 582854
rect 402102 582618 581546 582693
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 421008 579454
rect 421244 579218 555376 579454
rect 555612 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 421008 579134
rect 421244 578898 555376 579134
rect 555612 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 193210 547174
rect 193446 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 420328 547174
rect 420564 546938 556056 547174
rect 556292 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 193210 546854
rect 193446 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 420328 546854
rect 420564 546618 556056 546854
rect 556292 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 421008 543454
rect 421244 543218 555376 543454
rect 555612 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 421008 543134
rect 421244 542898 555376 543134
rect 555612 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 268706 522334
rect 268942 522098 269026 522334
rect 269262 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 268706 522014
rect 268942 521778 269026 522014
rect 269262 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 193210 511174
rect 193446 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 420328 511174
rect 420564 510938 556056 511174
rect 556292 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 193210 510854
rect 193446 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 420328 510854
rect 420564 510618 556056 510854
rect 556292 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 421008 507454
rect 421244 507218 555376 507454
rect 555612 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 421008 507134
rect 421244 506898 555376 507134
rect 555612 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 268706 486334
rect 268942 486098 269026 486334
rect 269262 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 268706 486014
rect 268942 485778 269026 486014
rect 269262 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 209610 439174
rect 209846 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 240330 439174
rect 240566 438938 271050 439174
rect 271286 438938 301770 439174
rect 302006 438938 332490 439174
rect 332726 438938 363210 439174
rect 363446 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 209610 438854
rect 209846 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 240330 438854
rect 240566 438618 271050 438854
rect 271286 438618 301770 438854
rect 302006 438618 332490 438854
rect 332726 438618 363210 438854
rect 363446 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 194250 435454
rect 194486 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 224970 435454
rect 225206 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 255690 435454
rect 255926 435218 286410 435454
rect 286646 435218 317130 435454
rect 317366 435218 347850 435454
rect 348086 435218 378570 435454
rect 378806 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 194250 435134
rect 194486 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 224970 435134
rect 225206 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 255690 435134
rect 255926 434898 286410 435134
rect 286646 434898 317130 435134
rect 317366 434898 347850 435134
rect 348086 434898 378570 435134
rect 378806 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 20328 403174
rect 20564 402938 156056 403174
rect 156292 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 209610 403174
rect 209846 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 240330 403174
rect 240566 402938 271050 403174
rect 271286 402938 301770 403174
rect 302006 402938 332490 403174
rect 332726 402938 363210 403174
rect 363446 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 420328 403174
rect 420564 402938 556056 403174
rect 556292 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 20328 402854
rect 20564 402618 156056 402854
rect 156292 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 209610 402854
rect 209846 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 240330 402854
rect 240566 402618 271050 402854
rect 271286 402618 301770 402854
rect 302006 402618 332490 402854
rect 332726 402618 363210 402854
rect 363446 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 420328 402854
rect 420564 402618 556056 402854
rect 556292 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 21008 399454
rect 21244 399218 155376 399454
rect 155612 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 194250 399454
rect 194486 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 224970 399454
rect 225206 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 255690 399454
rect 255926 399218 286410 399454
rect 286646 399218 317130 399454
rect 317366 399218 347850 399454
rect 348086 399218 378570 399454
rect 378806 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 421008 399454
rect 421244 399218 555376 399454
rect 555612 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 21008 399134
rect 21244 398898 155376 399134
rect 155612 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 194250 399134
rect 194486 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 224970 399134
rect 225206 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 255690 399134
rect 255926 398898 286410 399134
rect 286646 398898 317130 399134
rect 317366 398898 347850 399134
rect 348086 398898 378570 399134
rect 378806 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 421008 399134
rect 421244 398898 555376 399134
rect 555612 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 20328 367174
rect 20564 366938 156056 367174
rect 156292 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 209610 367174
rect 209846 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 240330 367174
rect 240566 366938 271050 367174
rect 271286 366938 301770 367174
rect 302006 366938 332490 367174
rect 332726 366938 363210 367174
rect 363446 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 420328 367174
rect 420564 366938 556056 367174
rect 556292 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 20328 366854
rect 20564 366618 156056 366854
rect 156292 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 209610 366854
rect 209846 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 240330 366854
rect 240566 366618 271050 366854
rect 271286 366618 301770 366854
rect 302006 366618 332490 366854
rect 332726 366618 363210 366854
rect 363446 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 420328 366854
rect 420564 366618 556056 366854
rect 556292 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 21008 363454
rect 21244 363218 155376 363454
rect 155612 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 194250 363454
rect 194486 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 224970 363454
rect 225206 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 255690 363454
rect 255926 363218 286410 363454
rect 286646 363218 317130 363454
rect 317366 363218 347850 363454
rect 348086 363218 378570 363454
rect 378806 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 421008 363454
rect 421244 363218 555376 363454
rect 555612 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 21008 363134
rect 21244 362898 155376 363134
rect 155612 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 194250 363134
rect 194486 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 224970 363134
rect 225206 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 255690 363134
rect 255926 362898 286410 363134
rect 286646 362898 317130 363134
rect 317366 362898 347850 363134
rect 348086 362898 378570 363134
rect 378806 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 421008 363134
rect 421244 362898 555376 363134
rect 555612 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 20328 331174
rect 20564 330938 156056 331174
rect 156292 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 209610 331174
rect 209846 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 240330 331174
rect 240566 330938 271050 331174
rect 271286 330938 301770 331174
rect 302006 330938 332490 331174
rect 332726 330938 363210 331174
rect 363446 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 420328 331174
rect 420564 330938 556056 331174
rect 556292 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 20328 330854
rect 20564 330618 156056 330854
rect 156292 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 209610 330854
rect 209846 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 240330 330854
rect 240566 330618 271050 330854
rect 271286 330618 301770 330854
rect 302006 330618 332490 330854
rect 332726 330618 363210 330854
rect 363446 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 420328 330854
rect 420564 330618 556056 330854
rect 556292 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 21008 327454
rect 21244 327218 155376 327454
rect 155612 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 194250 327454
rect 194486 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 224970 327454
rect 225206 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 255690 327454
rect 255926 327218 286410 327454
rect 286646 327218 317130 327454
rect 317366 327218 347850 327454
rect 348086 327218 378570 327454
rect 378806 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 421008 327454
rect 421244 327218 555376 327454
rect 555612 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 21008 327134
rect 21244 326898 155376 327134
rect 155612 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 194250 327134
rect 194486 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 224970 327134
rect 225206 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 255690 327134
rect 255926 326898 286410 327134
rect 286646 326898 317130 327134
rect 317366 326898 347850 327134
rect 348086 326898 378570 327134
rect 378806 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 421008 327134
rect 421244 326898 555376 327134
rect 555612 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 20328 295174
rect 20564 294938 156056 295174
rect 156292 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 209610 295174
rect 209846 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 240330 295174
rect 240566 294938 271050 295174
rect 271286 294938 301770 295174
rect 302006 294938 332490 295174
rect 332726 294938 363210 295174
rect 363446 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 420328 295174
rect 420564 294938 556056 295174
rect 556292 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 20328 294854
rect 20564 294618 156056 294854
rect 156292 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 209610 294854
rect 209846 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 240330 294854
rect 240566 294618 271050 294854
rect 271286 294618 301770 294854
rect 302006 294618 332490 294854
rect 332726 294618 363210 294854
rect 363446 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 420328 294854
rect 420564 294618 556056 294854
rect 556292 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 21008 291454
rect 21244 291218 155376 291454
rect 155612 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 194250 291454
rect 194486 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 224970 291454
rect 225206 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 255690 291454
rect 255926 291218 286410 291454
rect 286646 291218 317130 291454
rect 317366 291218 347850 291454
rect 348086 291218 378570 291454
rect 378806 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 421008 291454
rect 421244 291218 555376 291454
rect 555612 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 21008 291134
rect 21244 290898 155376 291134
rect 155612 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 194250 291134
rect 194486 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 224970 291134
rect 225206 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 255690 291134
rect 255926 290898 286410 291134
rect 286646 290898 317130 291134
rect 317366 290898 347850 291134
rect 348086 290898 378570 291134
rect 378806 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 421008 291134
rect 421244 290898 555376 291134
rect 555612 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 20328 259174
rect 20564 258938 156056 259174
rect 156292 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 209610 259174
rect 209846 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 240330 259174
rect 240566 258938 271050 259174
rect 271286 258938 301770 259174
rect 302006 258938 332490 259174
rect 332726 258938 363210 259174
rect 363446 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 420328 259174
rect 420564 258938 556056 259174
rect 556292 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 20328 258854
rect 20564 258618 156056 258854
rect 156292 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 209610 258854
rect 209846 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 240330 258854
rect 240566 258618 271050 258854
rect 271286 258618 301770 258854
rect 302006 258618 332490 258854
rect 332726 258618 363210 258854
rect 363446 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 420328 258854
rect 420564 258618 556056 258854
rect 556292 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 21008 255454
rect 21244 255218 155376 255454
rect 155612 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 194250 255454
rect 194486 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 224970 255454
rect 225206 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 255690 255454
rect 255926 255218 286410 255454
rect 286646 255218 317130 255454
rect 317366 255218 347850 255454
rect 348086 255218 378570 255454
rect 378806 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 421008 255454
rect 421244 255218 555376 255454
rect 555612 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 21008 255134
rect 21244 254898 155376 255134
rect 155612 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 194250 255134
rect 194486 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 224970 255134
rect 225206 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 255690 255134
rect 255926 254898 286410 255134
rect 286646 254898 317130 255134
rect 317366 254898 347850 255134
rect 348086 254898 378570 255134
rect 378806 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 421008 255134
rect 421244 254898 555376 255134
rect 555612 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 20328 223174
rect 20564 222938 156056 223174
rect 156292 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 420328 223174
rect 420564 222938 556056 223174
rect 556292 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 20328 222854
rect 20564 222618 156056 222854
rect 156292 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 420328 222854
rect 420564 222618 556056 222854
rect 556292 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 21008 219454
rect 21244 219218 155376 219454
rect 155612 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 421008 219454
rect 421244 219218 555376 219454
rect 555612 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 21008 219134
rect 21244 218898 155376 219134
rect 155612 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 421008 219134
rect 421244 218898 555376 219134
rect 555612 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 20328 187174
rect 20564 186938 156056 187174
rect 156292 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 420328 187174
rect 420564 186938 556056 187174
rect 556292 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 20328 186854
rect 20564 186618 156056 186854
rect 156292 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 420328 186854
rect 420564 186618 556056 186854
rect 556292 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 21008 183454
rect 21244 183218 155376 183454
rect 155612 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 421008 183454
rect 421244 183218 555376 183454
rect 555612 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 21008 183134
rect 21244 182898 155376 183134
rect 155612 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 421008 183134
rect 421244 182898 555376 183134
rect 555612 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 20328 151174
rect 20564 150938 156056 151174
rect 156292 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 420328 151174
rect 420564 150938 556056 151174
rect 556292 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 20328 150854
rect 20564 150618 156056 150854
rect 156292 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 420328 150854
rect 420564 150618 556056 150854
rect 556292 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 20328 115174
rect 20564 114938 156056 115174
rect 156292 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 420328 115174
rect 420564 114938 556056 115174
rect 556292 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 20328 114854
rect 20564 114618 156056 114854
rect 156292 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 420328 114854
rect 420564 114618 556056 114854
rect 556292 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 21008 111454
rect 21244 111218 155376 111454
rect 155612 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 421008 111454
rect 421244 111218 555376 111454
rect 555612 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 21008 111134
rect 21244 110898 155376 111134
rect 155612 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 421008 111134
rect 421244 110898 555376 111134
rect 555612 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 20328 79174
rect 20564 78938 156056 79174
rect 156292 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 420328 79174
rect 420564 78938 556056 79174
rect 556292 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 20328 78854
rect 20564 78618 156056 78854
rect 156292 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 420328 78854
rect 420564 78618 556056 78854
rect 556292 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 21008 75454
rect 21244 75218 155376 75454
rect 155612 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 421008 75454
rect 421244 75218 555376 75454
rect 555612 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 21008 75134
rect 21244 74898 155376 75134
rect 155612 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 421008 75134
rect 421244 74898 555376 75134
rect 555612 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use io_interface  IO_interface
timestamp 0
transform 1 0 190000 0 1 250000
box 1066 0 198850 200000
use sky130_sram_2kbyte_1rw1r_32x512_8  data_memory
timestamp 0
transform 1 0 420000 0 1 500000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory0
timestamp 0
transform 1 0 420000 0 1 150000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory1
timestamp 0
transform 1 0 420000 0 1 250000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory2
timestamp 0
transform 1 0 20000 0 1 150000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory3
timestamp 0
transform 1 0 20000 0 1 250000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory4
timestamp 0
transform 1 0 420000 0 1 50000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory5
timestamp 0
transform 1 0 420000 0 1 350000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory6
timestamp 0
transform 1 0 20000 0 1 50000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory7
timestamp 0
transform 1 0 20000 0 1 350000
box 0 0 136620 83308
use processor  uP
timestamp 0
transform 1 0 20000 0 1 500000
box 1066 0 178886 180000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 47940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 435244 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 47940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 435244 74414 501375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 678961 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 48064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 435244 110414 501375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 678961 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 48064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 435244 146414 501375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 678961 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 249743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 451537 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 249743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 451537 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 249743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 451537 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 48064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 435244 434414 498064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 585244 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 47940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 435244 470414 497940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 585244 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 47940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 435244 506414 497940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 585244 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 48064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 435244 542414 498064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 585244 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 47940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 435244 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 48064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 435244 81854 501375 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 678961 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 48064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 435244 117854 501375 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 678961 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 48064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 435244 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 250068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 449580 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 249743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 451537 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 249743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 451537 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 249743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 451537 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 47940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 435244 441854 497940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 585244 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 48064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 435244 477854 498064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 585244 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 47940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 435244 513854 497940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 585244 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 48064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 435244 549854 498064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 585244 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 48064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 435244 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 48064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 435244 89294 501375 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 48064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 435244 125294 501375 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 249743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 451537 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 249743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 451537 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 249743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 451537 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 47940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 435244 449294 497940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 585244 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 48064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 435244 485294 498064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 585244 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 47940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 435244 521294 497940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 585244 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 48064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 435244 557294 498064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 585244 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 48064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 435244 24734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 47940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 435244 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 48064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 435244 96734 501375 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 48064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 435244 132734 501375 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 250068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 449580 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 249743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 451537 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 249743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 451537 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 249743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 451537 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 48064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 435244 420734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 585244 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 47940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 435244 456734 497940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 585244 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 48064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 435244 492734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 585244 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 48064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 435244 528734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 585244 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 48064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 435244 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 47940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 435244 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 48064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 435244 93014 501375 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 48064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 435244 129014 501375 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 249743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 451537 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 249743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 451537 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 249743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 451537 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 47940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 435244 453014 497940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 585244 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 47940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 435244 489014 497940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 585244 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 48064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 435244 525014 498064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 585244 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 48064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 435244 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 47940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 435244 64454 501375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 48064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 435244 100454 501375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 48064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 435244 136454 501375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 249743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 451537 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 249743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 451537 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 249743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 451537 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 48064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 435244 424454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 585244 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 48064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 435244 460454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 585244 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 47940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 435244 496454 497940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 585244 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 48064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 435244 532454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 585244 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 47940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 435244 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 47940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 435244 78134 501375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 678961 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 47940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 435244 114134 501375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 678961 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 48064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 435244 150134 501375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 678961 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 451537 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 451537 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 451537 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 451537 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 48064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 435244 438134 498064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 585244 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 47940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 435244 474134 497940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 585244 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 48064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 435244 510134 498064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 585244 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 48064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 435244 546134 498064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 585244 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 48064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 435244 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 48064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 435244 85574 501375 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 678961 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 47940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 435244 121574 501375 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 678961 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 48064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 435244 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 500068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 679452 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 249743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 451537 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 249743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 451537 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 249743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 451537 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 47940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 435244 445574 497940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 585244 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 47940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 435244 481574 497940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 585244 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 48064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 435244 517574 498064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 585244 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 48064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 435244 553574 498064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 585244 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 155494 399336 155494 399336 0 vccd1
rlabel via4 189704 658776 189704 658776 0 vccd2
rlabel via4 197144 666216 197144 666216 0 vdda1
rlabel via4 168584 673656 168584 673656 0 vdda2
rlabel via4 164864 669936 164864 669936 0 vssa1
rlabel via4 172304 677376 172304 677376 0 vssa2
rlabel via4 156174 403056 156174 403056 0 vssd1
rlabel via4 157424 662496 157424 662496 0 vssd2
rlabel metal2 195024 679932 195024 679932 0 Serial_input
rlabel metal2 197218 679932 197218 679932 0 Serial_output
rlabel metal3 19719 58334 19719 58334 0 clk
rlabel metal4 436086 499818 436086 499818 0 data_mem_addr\[0\]
rlabel metal4 437174 499818 437174 499818 0 data_mem_addr\[1\]
rlabel metal2 296010 493816 296010 493816 0 data_mem_addr\[2\]
rlabel metal1 339894 461686 339894 461686 0 data_mem_addr\[3\]
rlabel metal1 273056 463250 273056 463250 0 data_mem_addr\[4\]
rlabel metal2 267950 462663 267950 462663 0 data_mem_addr\[5\]
rlabel metal2 269422 463377 269422 463377 0 data_mem_addr\[6\]
rlabel metal3 419735 535942 419735 535942 0 data_mem_addr\[7\]
rlabel metal1 279910 467194 279910 467194 0 data_mem_csb
rlabel metal4 448326 499818 448326 499818 0 data_read_data\[0\]
rlabel metal2 273509 449956 273509 449956 0 data_read_data\[10\]
rlabel metal2 274153 449956 274153 449956 0 data_read_data\[11\]
rlabel metal2 274981 449956 274981 449956 0 data_read_data\[12\]
rlabel metal2 275625 449956 275625 449956 0 data_read_data\[13\]
rlabel metal2 276407 449956 276407 449956 0 data_read_data\[14\]
rlabel metal2 277097 449956 277097 449956 0 data_read_data\[15\]
rlabel metal4 450774 499818 450774 499818 0 data_read_data\[1\]
rlabel metal1 358892 474062 358892 474062 0 data_read_data\[2\]
rlabel metal1 360548 475354 360548 475354 0 data_read_data\[3\]
rlabel metal1 362986 476782 362986 476782 0 data_read_data\[4\]
rlabel metal4 461110 499818 461110 499818 0 data_read_data\[5\]
rlabel metal4 463558 499818 463558 499818 0 data_read_data\[6\]
rlabel metal4 466006 499818 466006 499818 0 data_read_data\[7\]
rlabel metal4 468318 499818 468318 499818 0 data_read_data\[8\]
rlabel metal4 471038 499818 471038 499818 0 data_read_data\[9\]
rlabel metal4 438262 499818 438262 499818 0 data_wmask\[0\]
rlabel metal1 351256 483650 351256 483650 0 data_wmask\[1\]
rlabel metal1 352774 457470 352774 457470 0 data_wmask\[2\]
rlabel metal4 441798 499818 441798 499818 0 data_wmask\[3\]
rlabel metal4 443158 499818 443158 499818 0 data_write_data\[0\]
rlabel metal2 273785 449956 273785 449956 0 data_write_data\[10\]
rlabel metal2 274666 473032 274666 473032 0 data_write_data\[11\]
rlabel metal2 275257 449956 275257 449956 0 data_write_data\[12\]
rlabel metal2 276191 449956 276191 449956 0 data_write_data\[13\]
rlabel metal2 276729 449956 276729 449956 0 data_write_data\[14\]
rlabel metal2 277557 449956 277557 449956 0 data_write_data\[15\]
rlabel metal4 444246 499818 444246 499818 0 data_write_data\[1\]
rlabel metal4 445470 499818 445470 499818 0 data_write_data\[2\]
rlabel metal4 446558 499818 446558 499818 0 data_write_data\[3\]
rlabel metal4 447646 499818 447646 499818 0 data_write_data\[4\]
rlabel metal4 448734 499818 448734 499818 0 data_write_data\[5\]
rlabel metal4 450094 499818 450094 499818 0 data_write_data\[6\]
rlabel metal4 451076 498168 451076 498168 0 data_write_data\[7\]
rlabel metal1 361744 460258 361744 460258 0 data_write_data\[8\]
rlabel metal2 283590 475354 283590 475354 0 data_write_data\[9\]
rlabel metal2 277833 449956 277833 449956 0 dataw_enb
rlabel metal2 192632 679932 192632 679932 0 hlt
rlabel metal1 19596 249594 19596 249594 0 instr_mem_addr_9bit\[0\]
rlabel metal1 19504 249730 19504 249730 0 instr_mem_addr_9bit\[1\]
rlabel metal3 19719 78190 19719 78190 0 instr_mem_addr_9bit\[2\]
rlabel metal3 19719 79958 19719 79958 0 instr_mem_addr_9bit\[3\]
rlabel metal3 19719 81046 19719 81046 0 instr_mem_addr_9bit\[4\]
rlabel metal3 19903 82814 19903 82814 0 instr_mem_addr_9bit\[5\]
rlabel metal3 19719 83766 19719 83766 0 instr_mem_addr_9bit\[6\]
rlabel metal3 19719 385942 19719 385942 0 instr_mem_addr_9bit\[7\]
rlabel metal3 19719 386894 19719 386894 0 instr_mem_addr_9bit\[8\]
rlabel metal3 419735 158062 419735 158062 0 instr_mem_csb\[0\]
rlabel metal2 392702 356371 392702 356371 0 instr_mem_csb\[1\]
rlabel metal3 19811 158062 19811 158062 0 instr_mem_csb\[2\]
rlabel metal3 19719 258062 19719 258062 0 instr_mem_csb\[3\]
rlabel metal2 291962 451731 291962 451731 0 instr_mem_csb\[4\]
rlabel metal2 287546 451340 287546 451340 0 instr_mem_csb\[5\]
rlabel metal3 19903 58062 19903 58062 0 instr_mem_csb\[6\]
rlabel metal3 19903 358062 19903 358062 0 instr_mem_csb\[7\]
rlabel via3 448293 147628 448293 147628 0 instr_read_data0\[0\]
rlabel metal2 319095 449956 319095 449956 0 instr_read_data0\[10\]
rlabel metal2 322361 449956 322361 449956 0 instr_read_data0\[11\]
rlabel metal2 325818 450031 325818 450031 0 instr_read_data0\[12\]
rlabel metal2 328985 449956 328985 449956 0 instr_read_data0\[13\]
rlabel metal2 332297 449956 332297 449956 0 instr_read_data0\[14\]
rlabel metal2 412298 303382 412298 303382 0 instr_read_data0\[15\]
rlabel metal2 412482 303382 412482 303382 0 instr_read_data0\[16\]
rlabel metal2 412114 303110 412114 303110 0 instr_read_data0\[17\]
rlabel metal4 493478 149668 493478 149668 0 instr_read_data0\[18\]
rlabel metal2 412206 303042 412206 303042 0 instr_read_data0\[19\]
rlabel via3 450685 147628 450685 147628 0 instr_read_data0\[1\]
rlabel metal2 350842 450303 350842 450303 0 instr_read_data0\[20\]
rlabel metal2 353786 450167 353786 450167 0 instr_read_data0\[21\]
rlabel metal2 412390 303416 412390 303416 0 instr_read_data0\[22\]
rlabel metal2 412022 303212 412022 303212 0 instr_read_data0\[23\]
rlabel metal2 412574 299506 412574 299506 0 instr_read_data0\[24\]
rlabel metal2 365562 450218 365562 450218 0 instr_read_data0\[25\]
rlabel metal2 368605 449956 368605 449956 0 instr_read_data0\[26\]
rlabel metal2 371450 450116 371450 450116 0 instr_read_data0\[27\]
rlabel metal2 409630 299540 409630 299540 0 instr_read_data0\[28\]
rlabel metal2 409354 302430 409354 302430 0 instr_read_data0\[29\]
rlabel metal2 287769 449956 287769 449956 0 instr_read_data0\[2\]
rlabel metal2 406962 300645 406962 300645 0 instr_read_data0\[30\]
rlabel metal2 407054 299234 407054 299234 0 instr_read_data0\[31\]
rlabel metal2 292185 449956 292185 449956 0 instr_read_data0\[3\]
rlabel metal2 406502 302379 406502 302379 0 instr_read_data0\[4\]
rlabel metal2 406870 303416 406870 303416 0 instr_read_data0\[5\]
rlabel metal2 406778 301937 406778 301937 0 instr_read_data0\[6\]
rlabel metal2 406594 302668 406594 302668 0 instr_read_data0\[7\]
rlabel metal2 312425 449956 312425 449956 0 instr_read_data0\[8\]
rlabel metal2 315737 449956 315737 449956 0 instr_read_data0\[9\]
rlabel metal4 448326 249988 448326 249988 0 instr_read_data1\[0\]
rlabel metal2 319417 449956 319417 449956 0 instr_read_data1\[10\]
rlabel metal2 322874 450235 322874 450235 0 instr_read_data1\[11\]
rlabel metal2 326087 449956 326087 449956 0 instr_read_data1\[12\]
rlabel metal2 329353 449956 329353 449956 0 instr_read_data1\[13\]
rlabel metal2 332757 449956 332757 449956 0 instr_read_data1\[14\]
rlabel metal4 485998 249920 485998 249920 0 instr_read_data1\[15\]
rlabel metal4 488310 249920 488310 249920 0 instr_read_data1\[16\]
rlabel metal2 404110 353974 404110 353974 0 instr_read_data1\[17\]
rlabel metal2 404294 347820 404294 347820 0 instr_read_data1\[18\]
rlabel metal4 495926 249920 495926 249920 0 instr_read_data1\[19\]
rlabel metal4 450774 249988 450774 249988 0 instr_read_data1\[1\]
rlabel metal2 351065 449956 351065 449956 0 instr_read_data1\[20\]
rlabel metal2 354009 449956 354009 449956 0 instr_read_data1\[21\]
rlabel metal4 503542 249920 503542 249920 0 instr_read_data1\[22\]
rlabel metal4 505990 249852 505990 249852 0 instr_read_data1\[23\]
rlabel metal4 508574 249852 508574 249852 0 instr_read_data1\[24\]
rlabel metal2 365930 450252 365930 450252 0 instr_read_data1\[25\]
rlabel metal2 368874 450320 368874 450320 0 instr_read_data1\[26\]
rlabel metal2 371673 449956 371673 449956 0 instr_read_data1\[27\]
rlabel metal2 374617 449956 374617 449956 0 instr_read_data1\[28\]
rlabel metal4 520950 249852 520950 249852 0 instr_read_data1\[29\]
rlabel metal2 288137 449956 288137 449956 0 instr_read_data1\[2\]
rlabel metal4 523398 249988 523398 249988 0 instr_read_data1\[30\]
rlabel metal4 525982 249988 525982 249988 0 instr_read_data1\[31\]
rlabel metal4 456078 249852 456078 249852 0 instr_read_data1\[3\]
rlabel metal4 458526 249852 458526 249852 0 instr_read_data1\[4\]
rlabel metal4 461110 249852 461110 249852 0 instr_read_data1\[5\]
rlabel metal4 463558 249988 463558 249988 0 instr_read_data1\[6\]
rlabel metal4 466006 249988 466006 249988 0 instr_read_data1\[7\]
rlabel metal2 312793 449956 312793 449956 0 instr_read_data1\[8\]
rlabel metal2 405398 354688 405398 354688 0 instr_read_data1\[9\]
rlabel metal2 279673 449956 279673 449956 0 instr_read_data2\[0\]
rlabel metal2 319785 449956 319785 449956 0 instr_read_data2\[10\]
rlabel metal2 323189 449956 323189 449956 0 instr_read_data2\[11\]
rlabel metal2 326409 449956 326409 449956 0 instr_read_data2\[12\]
rlabel metal2 329919 449956 329919 449956 0 instr_read_data2\[13\]
rlabel metal2 333033 449956 333033 449956 0 instr_read_data2\[14\]
rlabel metal2 336345 449956 336345 449956 0 instr_read_data2\[15\]
rlabel metal2 339802 450150 339802 450150 0 instr_read_data2\[16\]
rlabel metal4 91030 149668 91030 149668 0 instr_read_data2\[17\]
rlabel metal4 93478 149804 93478 149804 0 instr_read_data2\[18\]
rlabel metal4 95926 149668 95926 149668 0 instr_read_data2\[19\]
rlabel metal2 284089 449956 284089 449956 0 instr_read_data2\[1\]
rlabel metal2 351578 450099 351578 450099 0 instr_read_data2\[20\]
rlabel metal2 354377 449956 354377 449956 0 instr_read_data2\[21\]
rlabel metal2 190946 347684 190946 347684 0 instr_read_data2\[22\]
rlabel metal2 156630 298469 156630 298469 0 instr_read_data2\[23\]
rlabel metal2 158194 301155 158194 301155 0 instr_read_data2\[24\]
rlabel metal2 366153 449956 366153 449956 0 instr_read_data2\[25\]
rlabel metal2 369097 449956 369097 449956 0 instr_read_data2\[26\]
rlabel metal2 372041 449956 372041 449956 0 instr_read_data2\[27\]
rlabel metal4 118502 149668 118502 149668 0 instr_read_data2\[28\]
rlabel metal4 120950 149804 120950 149804 0 instr_read_data2\[29\]
rlabel metal2 288551 449956 288551 449956 0 instr_read_data2\[2\]
rlabel metal4 123398 149668 123398 149668 0 instr_read_data2\[30\]
rlabel metal4 125982 149668 125982 149668 0 instr_read_data2\[31\]
rlabel metal4 56078 149804 56078 149804 0 instr_read_data2\[3\]
rlabel metal4 58526 149804 58526 149804 0 instr_read_data2\[4\]
rlabel metal2 180182 302345 180182 302345 0 instr_read_data2\[5\]
rlabel via3 63595 147628 63595 147628 0 instr_read_data2\[6\]
rlabel metal2 180090 302617 180090 302617 0 instr_read_data2\[7\]
rlabel metal2 313359 449956 313359 449956 0 instr_read_data2\[8\]
rlabel metal2 316473 449956 316473 449956 0 instr_read_data2\[9\]
rlabel metal2 180734 349928 180734 349928 0 instr_read_data3\[0\]
rlabel metal2 180550 352614 180550 352614 0 instr_read_data3\[10\]
rlabel metal4 76070 249988 76070 249988 0 instr_read_data3\[11\]
rlabel metal4 78518 249988 78518 249988 0 instr_read_data3\[12\]
rlabel metal4 80966 249988 80966 249988 0 instr_read_data3\[13\]
rlabel metal4 83550 249988 83550 249988 0 instr_read_data3\[14\]
rlabel metal2 177790 348279 177790 348279 0 instr_read_data3\[15\]
rlabel metal2 177606 353056 177606 353056 0 instr_read_data3\[16\]
rlabel metal2 177330 354824 177330 354824 0 instr_read_data3\[17\]
rlabel metal2 177698 354688 177698 354688 0 instr_read_data3\[18\]
rlabel metal4 95926 249920 95926 249920 0 instr_read_data3\[19\]
rlabel metal2 177974 349894 177974 349894 0 instr_read_data3\[1\]
rlabel metal4 98510 249920 98510 249920 0 instr_read_data3\[20\]
rlabel metal4 100958 249920 100958 249920 0 instr_read_data3\[21\]
rlabel metal2 174846 355470 174846 355470 0 instr_read_data3\[22\]
rlabel metal2 175214 354807 175214 354807 0 instr_read_data3\[23\]
rlabel metal2 174938 355504 174938 355504 0 instr_read_data3\[24\]
rlabel metal2 366521 449956 366521 449956 0 instr_read_data3\[25\]
rlabel metal4 113470 249852 113470 249852 0 instr_read_data3\[26\]
rlabel metal4 115918 249852 115918 249852 0 instr_read_data3\[27\]
rlabel metal4 118502 249988 118502 249988 0 instr_read_data3\[28\]
rlabel metal4 120950 249852 120950 249852 0 instr_read_data3\[29\]
rlabel metal2 288873 449956 288873 449956 0 instr_read_data3\[2\]
rlabel metal2 171810 355827 171810 355827 0 instr_read_data3\[30\]
rlabel metal2 389390 351169 389390 351169 0 instr_read_data3\[31\]
rlabel metal4 56078 249852 56078 249852 0 instr_read_data3\[3\]
rlabel metal4 58526 249852 58526 249852 0 instr_read_data3\[4\]
rlabel metal4 61110 249988 61110 249988 0 instr_read_data3\[5\]
rlabel metal4 63558 249988 63558 249988 0 instr_read_data3\[6\]
rlabel metal4 66006 249988 66006 249988 0 instr_read_data3\[7\]
rlabel metal2 313674 451459 313674 451459 0 instr_read_data3\[8\]
rlabel metal4 71038 249988 71038 249988 0 instr_read_data3\[9\]
rlabel metal2 405122 253555 405122 253555 0 instr_read_data4\[0\]
rlabel metal2 405214 250376 405214 250376 0 instr_read_data4\[10\]
rlabel metal2 405030 255323 405030 255323 0 instr_read_data4\[11\]
rlabel metal2 327237 449956 327237 449956 0 instr_read_data4\[12\]
rlabel metal2 330457 449956 330457 449956 0 instr_read_data4\[13\]
rlabel metal2 333769 449956 333769 449956 0 instr_read_data4\[14\]
rlabel metal2 407790 256173 407790 256173 0 instr_read_data4\[15\]
rlabel metal2 407974 255748 407974 255748 0 instr_read_data4\[16\]
rlabel metal2 410734 256309 410734 256309 0 instr_read_data4\[17\]
rlabel metal2 410642 256020 410642 256020 0 instr_read_data4\[18\]
rlabel metal2 407882 256428 407882 256428 0 instr_read_data4\[19\]
rlabel metal2 410550 255255 410550 255255 0 instr_read_data4\[1\]
rlabel metal2 352314 450915 352314 450915 0 instr_read_data4\[20\]
rlabel metal2 410826 256020 410826 256020 0 instr_read_data4\[21\]
rlabel metal4 503542 49892 503542 49892 0 instr_read_data4\[22\]
rlabel metal2 410918 252671 410918 252671 0 instr_read_data4\[23\]
rlabel metal4 508574 49824 508574 49824 0 instr_read_data4\[24\]
rlabel metal2 366889 449956 366889 449956 0 instr_read_data4\[25\]
rlabel metal2 369978 454094 369978 454094 0 instr_read_data4\[26\]
rlabel metal2 372823 449956 372823 449956 0 instr_read_data4\[27\]
rlabel metal2 375866 450847 375866 450847 0 instr_read_data4\[28\]
rlabel metal2 411930 249577 411930 249577 0 instr_read_data4\[29\]
rlabel metal2 289241 449956 289241 449956 0 instr_read_data4\[2\]
rlabel metal4 523398 50028 523398 50028 0 instr_read_data4\[30\]
rlabel metal4 525982 49824 525982 49824 0 instr_read_data4\[31\]
rlabel metal2 358754 450381 358754 450381 0 instr_read_data4\[3\]
rlabel metal1 357190 462366 357190 462366 0 instr_read_data4\[4\]
rlabel metal4 461110 50028 461110 50028 0 instr_read_data4\[5\]
rlabel metal2 403650 254524 403650 254524 0 instr_read_data4\[6\]
rlabel metal2 309166 461881 309166 461881 0 instr_read_data4\[7\]
rlabel metal2 313897 449956 313897 449956 0 instr_read_data4\[8\]
rlabel metal2 317209 449956 317209 449956 0 instr_read_data4\[9\]
rlabel metal4 448326 349968 448326 349968 0 instr_read_data5\[0\]
rlabel metal2 406226 405841 406226 405841 0 instr_read_data5\[10\]
rlabel metal4 476070 349968 476070 349968 0 instr_read_data5\[11\]
rlabel metal2 327658 451527 327658 451527 0 instr_read_data5\[12\]
rlabel metal4 480966 349968 480966 349968 0 instr_read_data5\[13\]
rlabel metal2 334183 449956 334183 449956 0 instr_read_data5\[14\]
rlabel metal4 485998 349968 485998 349968 0 instr_read_data5\[15\]
rlabel metal4 488310 349900 488310 349900 0 instr_read_data5\[16\]
rlabel metal4 491030 349900 491030 349900 0 instr_read_data5\[17\]
rlabel metal4 493478 349968 493478 349968 0 instr_read_data5\[18\]
rlabel metal1 389666 384982 389666 384982 0 instr_read_data5\[19\]
rlabel metal4 450774 349968 450774 349968 0 instr_read_data5\[1\]
rlabel metal2 352537 449956 352537 449956 0 instr_read_data5\[20\]
rlabel metal4 500958 349968 500958 349968 0 instr_read_data5\[21\]
rlabel metal4 503542 349968 503542 349968 0 instr_read_data5\[22\]
rlabel metal4 505990 349832 505990 349832 0 instr_read_data5\[23\]
rlabel metal2 364405 449956 364405 449956 0 instr_read_data5\[24\]
rlabel metal2 367402 451136 367402 451136 0 instr_read_data5\[25\]
rlabel metal2 370346 451306 370346 451306 0 instr_read_data5\[26\]
rlabel metal2 373290 450626 373290 450626 0 instr_read_data5\[27\]
rlabel metal2 392794 400214 392794 400214 0 instr_read_data5\[28\]
rlabel metal4 520950 349900 520950 349900 0 instr_read_data5\[29\]
rlabel metal2 289609 449956 289609 449956 0 instr_read_data5\[2\]
rlabel metal4 523398 349968 523398 349968 0 instr_read_data5\[30\]
rlabel metal4 525982 349968 525982 349968 0 instr_read_data5\[31\]
rlabel metal2 391230 400622 391230 400622 0 instr_read_data5\[3\]
rlabel metal4 458526 349968 458526 349968 0 instr_read_data5\[4\]
rlabel metal4 461110 349968 461110 349968 0 instr_read_data5\[5\]
rlabel metal4 463558 349832 463558 349832 0 instr_read_data5\[6\]
rlabel metal4 466006 349832 466006 349832 0 instr_read_data5\[7\]
rlabel metal2 314265 449956 314265 449956 0 instr_read_data5\[8\]
rlabel metal3 467820 347616 467820 347616 0 instr_read_data5\[9\]
rlabel metal2 281145 449956 281145 449956 0 instr_read_data6\[0\]
rlabel metal2 321257 449956 321257 449956 0 instr_read_data6\[10\]
rlabel metal4 76070 49878 76070 49878 0 instr_read_data6\[11\]
rlabel metal2 327881 449956 327881 449956 0 instr_read_data6\[12\]
rlabel metal2 331437 449956 331437 449956 0 instr_read_data6\[13\]
rlabel metal2 334505 449956 334505 449956 0 instr_read_data6\[14\]
rlabel metal2 337817 449956 337817 449956 0 instr_read_data6\[15\]
rlabel metal4 88310 49824 88310 49824 0 instr_read_data6\[16\]
rlabel metal4 91030 49892 91030 49892 0 instr_read_data6\[17\]
rlabel metal2 346610 462391 346610 462391 0 instr_read_data6\[18\]
rlabel metal4 95926 49892 95926 49892 0 instr_read_data6\[19\]
rlabel metal2 285805 449956 285805 449956 0 instr_read_data6\[1\]
rlabel metal2 352905 449956 352905 449956 0 instr_read_data6\[20\]
rlabel metal4 100958 50028 100958 50028 0 instr_read_data6\[21\]
rlabel metal2 358885 449956 358885 449956 0 instr_read_data6\[22\]
rlabel metal2 361737 449956 361737 449956 0 instr_read_data6\[23\]
rlabel metal2 364681 449956 364681 449956 0 instr_read_data6\[24\]
rlabel metal2 367625 449956 367625 449956 0 instr_read_data6\[25\]
rlabel metal2 370569 449956 370569 449956 0 instr_read_data6\[26\]
rlabel metal2 373513 449956 373513 449956 0 instr_read_data6\[27\]
rlabel metal4 118502 50028 118502 50028 0 instr_read_data6\[28\]
rlabel metal4 120950 49824 120950 49824 0 instr_read_data6\[29\]
rlabel metal2 290069 449956 290069 449956 0 instr_read_data6\[2\]
rlabel metal4 389252 248880 389252 248880 0 instr_read_data6\[30\]
rlabel metal2 388102 143493 388102 143493 0 instr_read_data6\[31\]
rlabel metal4 56078 49824 56078 49824 0 instr_read_data6\[3\]
rlabel metal4 58526 49824 58526 49824 0 instr_read_data6\[4\]
rlabel metal4 61110 50028 61110 50028 0 instr_read_data6\[5\]
rlabel metal4 63558 50028 63558 50028 0 instr_read_data6\[6\]
rlabel metal2 161138 255374 161138 255374 0 instr_read_data6\[7\]
rlabel metal2 314725 449956 314725 449956 0 instr_read_data6\[8\]
rlabel metal2 317945 449956 317945 449956 0 instr_read_data6\[9\]
rlabel metal2 191682 399245 191682 399245 0 instr_read_data7\[0\]
rlabel metal4 73622 349968 73622 349968 0 instr_read_data7\[10\]
rlabel metal4 76070 349832 76070 349832 0 instr_read_data7\[11\]
rlabel metal4 78518 349832 78518 349832 0 instr_read_data7\[12\]
rlabel metal4 80966 349968 80966 349968 0 instr_read_data7\[13\]
rlabel metal4 83550 349968 83550 349968 0 instr_read_data7\[14\]
rlabel metal2 177238 400758 177238 400758 0 instr_read_data7\[15\]
rlabel metal2 175122 401353 175122 401353 0 instr_read_data7\[16\]
rlabel metal2 172362 402016 172362 402016 0 instr_read_data7\[17\]
rlabel metal4 93478 349968 93478 349968 0 instr_read_data7\[18\]
rlabel metal4 95926 349832 95926 349832 0 instr_read_data7\[19\]
rlabel metal4 50774 349832 50774 349832 0 instr_read_data7\[1\]
rlabel metal4 98510 349968 98510 349968 0 instr_read_data7\[20\]
rlabel metal4 100958 349832 100958 349832 0 instr_read_data7\[21\]
rlabel metal4 103542 349968 103542 349968 0 instr_read_data7\[22\]
rlabel metal4 105990 349968 105990 349968 0 instr_read_data7\[23\]
rlabel metal2 365049 449956 365049 449956 0 instr_read_data7\[24\]
rlabel metal2 367993 449956 367993 449956 0 instr_read_data7\[25\]
rlabel metal4 113470 349968 113470 349968 0 instr_read_data7\[26\]
rlabel metal4 115918 349968 115918 349968 0 instr_read_data7\[27\]
rlabel metal4 118502 349968 118502 349968 0 instr_read_data7\[28\]
rlabel metal4 120950 349968 120950 349968 0 instr_read_data7\[29\]
rlabel metal2 190946 348449 190946 348449 0 instr_read_data7\[2\]
rlabel metal2 156722 403240 156722 403240 0 instr_read_data7\[30\]
rlabel metal2 159850 403308 159850 403308 0 instr_read_data7\[31\]
rlabel metal4 56078 349832 56078 349832 0 instr_read_data7\[3\]
rlabel metal4 58526 349832 58526 349832 0 instr_read_data7\[4\]
rlabel metal2 158562 400299 158562 400299 0 instr_read_data7\[5\]
rlabel metal2 165370 397936 165370 397936 0 instr_read_data7\[6\]
rlabel metal2 165094 401132 165094 401132 0 instr_read_data7\[7\]
rlabel metal2 157918 400265 157918 400265 0 instr_read_data7\[8\]
rlabel metal2 190670 347276 190670 347276 0 instr_read_data7\[9\]
rlabel metal4 38262 249988 38262 249988 0 instr_wmask\[0\]
rlabel metal3 18791 249764 18791 249764 0 instr_wmask\[1\]
rlabel metal4 40574 249988 40574 249988 0 instr_wmask\[2\]
rlabel metal4 41798 249988 41798 249988 0 instr_wmask\[3\]
rlabel metal4 43158 249988 43158 249988 0 instr_write_data\[0\]
rlabel via1 55246 346715 55246 346715 0 instr_write_data\[10\]
rlabel metal4 55942 249988 55942 249988 0 instr_write_data\[11\]
rlabel metal1 19182 234974 19182 234974 0 instr_write_data\[12\]
rlabel metal4 58118 249988 58118 249988 0 instr_write_data\[13\]
rlabel metal4 59478 249988 59478 249988 0 instr_write_data\[14\]
rlabel metal4 60702 249988 60702 249988 0 instr_write_data\[15\]
rlabel metal4 44246 249988 44246 249988 0 instr_write_data\[1\]
rlabel metal4 45470 249988 45470 249988 0 instr_write_data\[2\]
rlabel metal4 446558 249988 446558 249988 0 instr_write_data\[3\]
rlabel metal4 447646 249988 447646 249988 0 instr_write_data\[4\]
rlabel metal4 448734 249988 448734 249988 0 instr_write_data\[5\]
rlabel metal4 450094 249988 450094 249988 0 instr_write_data\[6\]
rlabel metal1 18492 235110 18492 235110 0 instr_write_data\[7\]
rlabel metal2 190854 348585 190854 348585 0 instr_write_data\[8\]
rlabel metal2 190946 400452 190946 400452 0 instr_write_data\[9\]
rlabel metal3 19719 59966 19719 59966 0 instrw_enb
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel via2 580198 458133 580198 458133 0 io_in[10]
rlabel metal2 558302 504730 558302 504730 0 io_in[11]
rlabel metal2 580198 563703 580198 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel metal2 231150 567562 231150 567562 0 io_in[14]
rlabel metal1 558946 699686 558946 699686 0 io_in[15]
rlabel metal1 352682 584426 352682 584426 0 io_in[16]
rlabel metal2 211830 460920 211830 460920 0 io_in[17]
rlabel metal2 364366 602691 364366 602691 0 io_in[18]
rlabel metal2 214314 460920 214314 460920 0 io_in[19]
rlabel metal2 194810 451187 194810 451187 0 io_in[1]
rlabel metal2 215641 449956 215641 449956 0 io_in[20]
rlabel metal2 216791 449956 216791 449956 0 io_in[21]
rlabel metal2 217849 449956 217849 449956 0 io_in[22]
rlabel metal2 218953 449956 218953 449956 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 1556 632060 1556 632060 0 io_in[25]
rlabel metal3 1832 579972 1832 579972 0 io_in[26]
rlabel metal3 1648 527884 1648 527884 0 io_in[27]
rlabel metal3 1878 475660 1878 475660 0 io_in[28]
rlabel metal3 1786 423572 1786 423572 0 io_in[29]
rlabel metal2 195914 451051 195914 451051 0 io_in[2]
rlabel metal3 2154 371348 2154 371348 0 io_in[30]
rlabel metal2 193154 449735 193154 449735 0 io_in[31]
rlabel metal3 1970 267172 1970 267172 0 io_in[32]
rlabel metal3 1832 214948 1832 214948 0 io_in[33]
rlabel metal2 231097 449956 231097 449956 0 io_in[34]
rlabel metal3 1740 110636 1740 110636 0 io_in[35]
rlabel metal2 233397 449956 233397 449956 0 io_in[36]
rlabel metal2 234409 449956 234409 449956 0 io_in[37]
rlabel metal3 582230 126004 582230 126004 0 io_in[3]
rlabel metal3 582046 165852 582046 165852 0 io_in[4]
rlabel metal3 582000 205700 582000 205700 0 io_in[5]
rlabel metal3 582046 245548 582046 245548 0 io_in[6]
rlabel metal3 581862 298724 581862 298724 0 io_in[7]
rlabel metal2 580106 352563 580106 352563 0 io_in[8]
rlabel metal2 580106 405297 580106 405297 0 io_in[9]
rlabel metal3 193959 449276 193959 449276 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 563730 505410 563730 505410 0 io_oeb[11]
rlabel metal2 579830 590835 579830 590835 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 527206 701940 527206 701940 0 io_oeb[15]
rlabel metal2 462346 645364 462346 645364 0 io_oeb[16]
rlabel metal1 304750 501602 304750 501602 0 io_oeb[17]
rlabel metal1 331890 703018 331890 703018 0 io_oeb[18]
rlabel metal1 267030 697578 267030 697578 0 io_oeb[19]
rlabel metal2 308614 249917 308614 249917 0 io_oeb[1]
rlabel metal2 216009 449956 216009 449956 0 io_oeb[20]
rlabel metal2 217113 449956 217113 449956 0 io_oeb[21]
rlabel metal2 218217 449956 218217 449956 0 io_oeb[22]
rlabel metal1 9246 699686 9246 699686 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 1786 606084 1786 606084 0 io_oeb[25]
rlabel metal3 1832 553860 1832 553860 0 io_oeb[26]
rlabel metal3 1832 501772 1832 501772 0 io_oeb[27]
rlabel metal3 1924 449548 1924 449548 0 io_oeb[28]
rlabel metal3 2200 397460 2200 397460 0 io_oeb[29]
rlabel metal3 581908 112812 581908 112812 0 io_oeb[2]
rlabel metal2 191866 397681 191866 397681 0 io_oeb[30]
rlabel metal3 2016 293148 2016 293148 0 io_oeb[31]
rlabel metal2 229257 449956 229257 449956 0 io_oeb[32]
rlabel metal2 230559 449956 230559 449956 0 io_oeb[33]
rlabel metal3 1924 136748 1924 136748 0 io_oeb[34]
rlabel metal2 232569 449956 232569 449956 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal3 581954 152660 581954 152660 0 io_oeb[3]
rlabel metal1 578726 193154 578726 193154 0 io_oeb[4]
rlabel metal1 578818 233206 578818 233206 0 io_oeb[5]
rlabel metal3 582184 272204 582184 272204 0 io_oeb[6]
rlabel metal2 563730 393346 563730 393346 0 io_oeb[7]
rlabel metal2 580106 378947 580106 378947 0 io_oeb[8]
rlabel metal2 580106 431749 580106 431749 0 io_oeb[9]
rlabel metal3 194097 450364 194097 450364 0 io_out[0]
rlabel metal2 580014 471019 580014 471019 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal3 581908 577660 581908 577660 0 io_out[12]
rlabel metal2 580198 630751 580198 630751 0 io_out[13]
rlabel metal2 580198 683519 580198 683519 0 io_out[14]
rlabel metal2 542386 645497 542386 645497 0 io_out[15]
rlabel metal2 371910 603058 371910 603058 0 io_out[16]
rlabel metal1 313122 700298 313122 700298 0 io_out[17]
rlabel metal1 347254 699686 347254 699686 0 io_out[18]
rlabel metal2 215418 470992 215418 470992 0 io_out[19]
rlabel metal2 193246 449599 193246 449599 0 io_out[1]
rlabel metal2 216377 449956 216377 449956 0 io_out[20]
rlabel metal2 217481 449956 217481 449956 0 io_out[21]
rlabel metal2 218585 449956 218585 449956 0 io_out[22]
rlabel metal2 23828 703596 23828 703596 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal3 1924 514828 1924 514828 0 io_out[27]
rlabel metal3 1786 462604 1786 462604 0 io_out[28]
rlabel metal3 1832 410516 1832 410516 0 io_out[29]
rlabel metal1 578634 100674 578634 100674 0 io_out[2]
rlabel metal3 1878 358428 1878 358428 0 io_out[30]
rlabel metal3 2062 306204 2062 306204 0 io_out[31]
rlabel metal3 1924 254116 1924 254116 0 io_out[32]
rlabel metal2 230775 449956 230775 449956 0 io_out[33]
rlabel metal2 231925 449956 231925 449956 0 io_out[34]
rlabel metal3 1924 97580 1924 97580 0 io_out[35]
rlabel metal3 1878 58548 1878 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel metal1 578634 139366 578634 139366 0 io_out[3]
rlabel metal1 578910 179350 578910 179350 0 io_out[4]
rlabel metal1 578956 219198 578956 219198 0 io_out[5]
rlabel metal3 582092 258876 582092 258876 0 io_out[6]
rlabel metal3 581770 312052 581770 312052 0 io_out[7]
rlabel metal3 582138 365092 582138 365092 0 io_out[8]
rlabel metal2 559590 440334 559590 440334 0 io_out[9]
rlabel metal2 194665 250036 194665 250036 0 la_data_in[0]
rlabel metal2 197478 146040 197478 146040 0 la_data_out[0]
rlabel metal2 481758 3968 481758 3968 0 la_data_out[100]
rlabel metal2 485254 1622 485254 1622 0 la_data_out[101]
rlabel metal2 488842 4648 488842 4648 0 la_data_out[102]
rlabel metal2 339565 250036 339565 250036 0 la_data_out[103]
rlabel metal2 340945 250036 340945 250036 0 la_data_out[104]
rlabel metal2 342325 250036 342325 250036 0 la_data_out[105]
rlabel metal2 502688 16560 502688 16560 0 la_data_out[106]
rlabel metal2 345085 250036 345085 250036 0 la_data_out[107]
rlabel metal2 346465 250036 346465 250036 0 la_data_out[108]
rlabel metal2 347845 250036 347845 250036 0 la_data_out[109]
rlabel metal2 211225 250036 211225 250036 0 la_data_out[10]
rlabel metal2 349225 250036 349225 250036 0 la_data_out[110]
rlabel metal2 350605 250036 350605 250036 0 la_data_out[111]
rlabel metal2 351985 250036 351985 250036 0 la_data_out[112]
rlabel metal2 353365 250036 353365 250036 0 la_data_out[113]
rlabel metal2 354745 250036 354745 250036 0 la_data_out[114]
rlabel metal2 356125 250036 356125 250036 0 la_data_out[115]
rlabel metal2 538430 2642 538430 2642 0 la_data_out[116]
rlabel metal2 542018 2608 542018 2608 0 la_data_out[117]
rlabel metal2 545514 2574 545514 2574 0 la_data_out[118]
rlabel metal2 361645 250036 361645 250036 0 la_data_out[119]
rlabel metal2 212658 247496 212658 247496 0 la_data_out[11]
rlabel metal2 363025 250036 363025 250036 0 la_data_out[120]
rlabel metal2 364405 250036 364405 250036 0 la_data_out[121]
rlabel metal2 559774 1622 559774 1622 0 la_data_out[122]
rlabel metal2 367165 250036 367165 250036 0 la_data_out[123]
rlabel metal2 368545 250036 368545 250036 0 la_data_out[124]
rlabel metal2 369925 250036 369925 250036 0 la_data_out[125]
rlabel metal2 371305 250036 371305 250036 0 la_data_out[126]
rlabel metal2 577438 2234 577438 2234 0 la_data_out[127]
rlabel metal2 213985 250036 213985 250036 0 la_data_out[12]
rlabel metal2 172953 340 172953 340 0 la_data_out[13]
rlabel metal2 216745 250036 216745 250036 0 la_data_out[14]
rlabel metal2 218125 250036 218125 250036 0 la_data_out[15]
rlabel metal2 219505 250036 219505 250036 0 la_data_out[16]
rlabel metal2 187121 340 187121 340 0 la_data_out[17]
rlabel metal2 190663 340 190663 340 0 la_data_out[18]
rlabel metal2 194442 2608 194442 2608 0 la_data_out[19]
rlabel metal2 198805 250036 198805 250036 0 la_data_out[1]
rlabel metal2 197662 16560 197662 16560 0 la_data_out[20]
rlabel metal2 226405 250036 226405 250036 0 la_data_out[21]
rlabel metal2 218730 125562 218730 125562 0 la_data_out[22]
rlabel metal2 229218 248924 229218 248924 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215694 1962 215694 1962 0 la_data_out[25]
rlabel metal2 219282 1996 219282 1996 0 la_data_out[26]
rlabel metal2 234685 250036 234685 250036 0 la_data_out[27]
rlabel metal2 236118 248856 236118 248856 0 la_data_out[28]
rlabel metal2 229862 1928 229862 1928 0 la_data_out[29]
rlabel metal2 134037 340 134037 340 0 la_data_out[2]
rlabel metal2 233450 1792 233450 1792 0 la_data_out[30]
rlabel metal2 237038 1690 237038 1690 0 la_data_out[31]
rlabel metal2 240534 1928 240534 1928 0 la_data_out[32]
rlabel metal2 244122 1928 244122 1928 0 la_data_out[33]
rlabel metal2 247618 1962 247618 1962 0 la_data_out[34]
rlabel metal2 251206 1928 251206 1928 0 la_data_out[35]
rlabel metal2 254702 1894 254702 1894 0 la_data_out[36]
rlabel metal2 248485 250036 248485 250036 0 la_data_out[37]
rlabel metal2 249865 250036 249865 250036 0 la_data_out[38]
rlabel metal2 251245 250036 251245 250036 0 la_data_out[39]
rlabel metal2 137678 1894 137678 1894 0 la_data_out[3]
rlabel metal2 252625 250036 252625 250036 0 la_data_out[40]
rlabel metal2 254005 250036 254005 250036 0 la_data_out[41]
rlabel metal2 255385 250036 255385 250036 0 la_data_out[42]
rlabel metal2 256765 250036 256765 250036 0 la_data_out[43]
rlabel metal2 258145 250036 258145 250036 0 la_data_out[44]
rlabel metal2 259525 250036 259525 250036 0 la_data_out[45]
rlabel metal2 290214 1928 290214 1928 0 la_data_out[46]
rlabel metal2 293710 1690 293710 1690 0 la_data_out[47]
rlabel metal2 294078 5270 294078 5270 0 la_data_out[48]
rlabel metal2 265045 250036 265045 250036 0 la_data_out[49]
rlabel metal2 141266 1928 141266 1928 0 la_data_out[4]
rlabel metal2 266425 250036 266425 250036 0 la_data_out[50]
rlabel metal2 267805 250036 267805 250036 0 la_data_out[51]
rlabel metal2 269185 250036 269185 250036 0 la_data_out[52]
rlabel metal2 270565 250036 270565 250036 0 la_data_out[53]
rlabel metal1 272964 247078 272964 247078 0 la_data_out[54]
rlabel metal2 273325 250036 273325 250036 0 la_data_out[55]
rlabel metal2 274705 250036 274705 250036 0 la_data_out[56]
rlabel metal2 276085 250036 276085 250036 0 la_data_out[57]
rlabel metal2 332718 3968 332718 3968 0 la_data_out[58]
rlabel metal2 278845 250036 278845 250036 0 la_data_out[59]
rlabel metal2 144762 1962 144762 1962 0 la_data_out[5]
rlabel metal2 280225 250036 280225 250036 0 la_data_out[60]
rlabel metal2 281605 250036 281605 250036 0 la_data_out[61]
rlabel metal2 346978 2676 346978 2676 0 la_data_out[62]
rlabel metal2 350474 2642 350474 2642 0 la_data_out[63]
rlabel metal2 354062 2608 354062 2608 0 la_data_out[64]
rlabel metal2 287125 250036 287125 250036 0 la_data_out[65]
rlabel metal2 288505 250036 288505 250036 0 la_data_out[66]
rlabel metal2 289938 248550 289938 248550 0 la_data_out[67]
rlabel metal2 291265 250036 291265 250036 0 la_data_out[68]
rlabel metal2 292645 250036 292645 250036 0 la_data_out[69]
rlabel metal2 148350 1996 148350 1996 0 la_data_out[6]
rlabel metal2 294025 250036 294025 250036 0 la_data_out[70]
rlabel metal2 295405 250036 295405 250036 0 la_data_out[71]
rlabel metal2 296785 250036 296785 250036 0 la_data_out[72]
rlabel metal2 385986 2166 385986 2166 0 la_data_out[73]
rlabel metal2 389344 16560 389344 16560 0 la_data_out[74]
rlabel metal2 393070 3356 393070 3356 0 la_data_out[75]
rlabel metal2 302305 250036 302305 250036 0 la_data_out[76]
rlabel metal2 303685 250036 303685 250036 0 la_data_out[77]
rlabel metal2 403650 2132 403650 2132 0 la_data_out[78]
rlabel metal2 306498 248924 306498 248924 0 la_data_out[79]
rlabel metal2 151846 2030 151846 2030 0 la_data_out[7]
rlabel metal2 307878 248890 307878 248890 0 la_data_out[80]
rlabel metal2 309258 248856 309258 248856 0 la_data_out[81]
rlabel metal2 310585 250036 310585 250036 0 la_data_out[82]
rlabel metal1 312984 247078 312984 247078 0 la_data_out[83]
rlabel metal2 313345 250036 313345 250036 0 la_data_out[84]
rlabel metal2 314725 250036 314725 250036 0 la_data_out[85]
rlabel metal2 316105 250036 316105 250036 0 la_data_out[86]
rlabel metal2 317485 250036 317485 250036 0 la_data_out[87]
rlabel metal2 318865 250036 318865 250036 0 la_data_out[88]
rlabel metal2 442152 16560 442152 16560 0 la_data_out[89]
rlabel metal2 155434 2064 155434 2064 0 la_data_out[8]
rlabel metal2 446009 340 446009 340 0 la_data_out[90]
rlabel metal2 449834 1554 449834 1554 0 la_data_out[91]
rlabel metal2 324385 250036 324385 250036 0 la_data_out[92]
rlabel metal1 327474 247078 327474 247078 0 la_data_out[93]
rlabel metal2 327145 250036 327145 250036 0 la_data_out[94]
rlabel metal2 328525 250036 328525 250036 0 la_data_out[95]
rlabel metal2 329905 250036 329905 250036 0 la_data_out[96]
rlabel metal2 331285 250036 331285 250036 0 la_data_out[97]
rlabel metal2 332718 248550 332718 248550 0 la_data_out[98]
rlabel metal2 334045 250036 334045 250036 0 la_data_out[99]
rlabel metal2 158930 2098 158930 2098 0 la_data_out[9]
rlabel metal1 195684 247078 195684 247078 0 la_oenb[0]
rlabel metal3 156588 229224 156588 229224 0 low
rlabel metal2 154760 500140 154760 500140 0 reset
rlabel metal2 389206 463539 389206 463539 0 start
rlabel metal2 92168 679932 92168 679932 0 uP_data_mem_addr\[0\]
rlabel metal2 94560 679932 94560 679932 0 uP_data_mem_addr\[1\]
rlabel metal2 96952 679932 96952 679932 0 uP_data_mem_addr\[2\]
rlabel metal2 99252 679932 99252 679932 0 uP_data_mem_addr\[3\]
rlabel metal2 101736 679932 101736 679932 0 uP_data_mem_addr\[4\]
rlabel metal2 104128 679932 104128 679932 0 uP_data_mem_addr\[5\]
rlabel metal2 106520 679932 106520 679932 0 uP_data_mem_addr\[6\]
rlabel metal2 248761 449956 248761 449956 0 uP_data_mem_addr\[7\]
rlabel via1 187818 679405 187818 679405 0 uP_dataw_en
rlabel metal2 22372 679252 22372 679252 0 uP_instr\[0\]
rlabel metal2 253545 449956 253545 449956 0 uP_instr\[10\]
rlabel metal2 75424 679932 75424 679932 0 uP_instr\[11\]
rlabel metal2 80010 679932 80010 679932 0 uP_instr\[12\]
rlabel metal2 137310 681224 137310 681224 0 uP_instr\[13\]
rlabel metal2 98670 680680 98670 680680 0 uP_instr\[14\]
rlabel metal1 93840 679218 93840 679218 0 uP_instr\[15\]
rlabel metal2 79074 680663 79074 680663 0 uP_instr\[1\]
rlabel metal2 32368 679932 32368 679932 0 uP_instr\[2\]
rlabel metal2 37106 679932 37106 679932 0 uP_instr\[3\]
rlabel metal2 41936 679932 41936 679932 0 uP_instr\[4\]
rlabel metal2 46720 679932 46720 679932 0 uP_instr\[5\]
rlabel metal2 51504 679932 51504 679932 0 uP_instr\[6\]
rlabel metal2 56288 679932 56288 679932 0 uP_instr\[7\]
rlabel metal2 61072 679932 61072 679932 0 uP_instr\[8\]
rlabel metal2 100786 681632 100786 681632 0 uP_instr\[9\]
rlabel metal2 25192 679932 25192 679932 0 uP_instr_mem_addr\[0\]
rlabel metal2 72986 679932 72986 679932 0 uP_instr_mem_addr\[10\]
rlabel metal2 77816 679932 77816 679932 0 uP_instr_mem_addr\[11\]
rlabel metal2 82600 679932 82600 679932 0 uP_instr_mem_addr\[12\]
rlabel metal2 29976 679932 29976 679932 0 uP_instr_mem_addr\[1\]
rlabel metal2 34760 679932 34760 679932 0 uP_instr_mem_addr\[2\]
rlabel metal2 39544 679932 39544 679932 0 uP_instr_mem_addr\[3\]
rlabel metal2 44130 679932 44130 679932 0 uP_instr_mem_addr\[4\]
rlabel metal2 49112 679932 49112 679932 0 uP_instr_mem_addr\[5\]
rlabel metal2 53698 679796 53698 679796 0 uP_instr_mem_addr\[6\]
rlabel metal2 58680 679932 58680 679932 0 uP_instr_mem_addr\[7\]
rlabel metal2 63372 679932 63372 679932 0 uP_instr_mem_addr\[8\]
rlabel metal2 252731 449820 252731 449820 0 uP_instr_mem_addr\[9\]
rlabel metal2 111304 679932 111304 679932 0 uP_read_data\[0\]
rlabel via1 135194 679405 135194 679405 0 uP_read_data\[10\]
rlabel metal2 137616 679932 137616 679932 0 uP_read_data\[11\]
rlabel metal2 140008 679932 140008 679932 0 uP_read_data\[12\]
rlabel metal2 142400 679932 142400 679932 0 uP_read_data\[13\]
rlabel metal2 144746 679932 144746 679932 0 uP_read_data\[14\]
rlabel metal2 147184 679932 147184 679932 0 uP_read_data\[15\]
rlabel metal1 113850 679252 113850 679252 0 uP_read_data\[1\]
rlabel metal1 116058 679286 116058 679286 0 uP_read_data\[2\]
rlabel metal2 118480 679932 118480 679932 0 uP_read_data\[3\]
rlabel via1 121026 679405 121026 679405 0 uP_read_data\[4\]
rlabel metal2 123264 679932 123264 679932 0 uP_read_data\[5\]
rlabel metal2 125458 679796 125458 679796 0 uP_read_data\[6\]
rlabel metal2 249957 449956 249957 449956 0 uP_read_data\[7\]
rlabel metal2 251429 449956 251429 449956 0 uP_read_data\[8\]
rlabel metal2 132832 679932 132832 679932 0 uP_read_data\[9\]
rlabel metal2 149576 679932 149576 679932 0 uP_write_data\[0\]
rlabel metal2 173496 679932 173496 679932 0 uP_write_data\[10\]
rlabel metal2 175888 679932 175888 679932 0 uP_write_data\[11\]
rlabel metal2 178280 679932 178280 679932 0 uP_write_data\[12\]
rlabel metal2 180580 679932 180580 679932 0 uP_write_data\[13\]
rlabel metal2 183064 679932 183064 679932 0 uP_write_data\[14\]
rlabel metal2 185456 679932 185456 679932 0 uP_write_data\[15\]
rlabel via1 151938 679405 151938 679405 0 uP_write_data\[1\]
rlabel metal2 154268 679932 154268 679932 0 uP_write_data\[2\]
rlabel metal2 156752 679932 156752 679932 0 uP_write_data\[3\]
rlabel metal2 159144 679932 159144 679932 0 uP_write_data\[4\]
rlabel metal2 161368 680075 161368 680075 0 uP_write_data\[5\]
rlabel metal2 248485 449956 248485 449956 0 uP_write_data\[6\]
rlabel metal2 250233 449956 250233 449956 0 uP_write_data\[7\]
rlabel metal2 251705 449956 251705 449956 0 uP_write_data\[8\]
rlabel metal2 253177 449956 253177 449956 0 uP_write_data\[9\]
rlabel metal2 581026 1894 581026 1894 0 user_irq[0]
rlabel metal2 582222 1792 582222 1792 0 user_irq[1]
rlabel metal2 582912 16560 582912 16560 0 user_irq[2]
rlabel metal2 598 2234 598 2234 0 wb_clk_i
rlabel metal2 1702 1928 1702 1928 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
