magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< metal1 >>
rect 1465 2168 1471 2220
rect 1523 2168 1529 2220
rect 1570 1130 1604 2256
rect 1646 1142 1674 2256
rect 2713 2168 2719 2220
rect 2771 2168 2777 2220
rect 1793 2016 1799 2068
rect 1851 2016 1857 2068
rect 1711 1242 1717 1294
rect 1769 1242 1775 1294
rect 2818 1130 2852 2256
rect 2894 1142 2922 2256
rect 3961 2168 3967 2220
rect 4019 2168 4025 2220
rect 3041 2016 3047 2068
rect 3099 2016 3105 2068
rect 2959 1242 2965 1294
rect 3017 1242 3023 1294
rect 4066 1130 4100 2256
rect 4142 1142 4170 2256
rect 5209 2168 5215 2220
rect 5267 2168 5273 2220
rect 4289 2016 4295 2068
rect 4347 2016 4353 2068
rect 4207 1242 4213 1294
rect 4265 1242 4271 1294
rect 5314 1130 5348 2256
rect 5390 1142 5418 2256
rect 6457 2168 6463 2220
rect 6515 2168 6521 2220
rect 5537 2016 5543 2068
rect 5595 2016 5601 2068
rect 5455 1242 5461 1294
rect 5513 1242 5519 1294
rect 6562 1130 6596 2256
rect 6638 1142 6666 2256
rect 7705 2168 7711 2220
rect 7763 2168 7769 2220
rect 6785 2016 6791 2068
rect 6843 2016 6849 2068
rect 6703 1242 6709 1294
rect 6761 1242 6767 1294
rect 7810 1130 7844 2256
rect 7886 1142 7914 2256
rect 8953 2168 8959 2220
rect 9011 2168 9017 2220
rect 8033 2016 8039 2068
rect 8091 2016 8097 2068
rect 7951 1242 7957 1294
rect 8009 1242 8015 1294
rect 9058 1130 9092 2256
rect 9134 1142 9162 2256
rect 10201 2168 10207 2220
rect 10259 2168 10265 2220
rect 9281 2016 9287 2068
rect 9339 2016 9345 2068
rect 9199 1242 9205 1294
rect 9257 1242 9263 1294
rect 10306 1130 10340 2256
rect 10382 1142 10410 2256
rect 11449 2168 11455 2220
rect 11507 2168 11513 2220
rect 10529 2016 10535 2068
rect 10587 2016 10593 2068
rect 10447 1242 10453 1294
rect 10505 1242 10511 1294
rect 11554 1130 11588 2256
rect 11630 1142 11658 2256
rect 12697 2168 12703 2220
rect 12755 2168 12761 2220
rect 11777 2016 11783 2068
rect 11835 2016 11841 2068
rect 11695 1242 11701 1294
rect 11753 1242 11759 1294
rect 12802 1130 12836 2256
rect 12878 1142 12906 2256
rect 13945 2168 13951 2220
rect 14003 2168 14009 2220
rect 13025 2016 13031 2068
rect 13083 2016 13089 2068
rect 12943 1242 12949 1294
rect 13001 1242 13007 1294
rect 14050 1130 14084 2256
rect 14126 1142 14154 2256
rect 15193 2168 15199 2220
rect 15251 2168 15257 2220
rect 14273 2016 14279 2068
rect 14331 2016 14337 2068
rect 14191 1242 14197 1294
rect 14249 1242 14255 1294
rect 15298 1130 15332 2256
rect 15374 1142 15402 2256
rect 16441 2168 16447 2220
rect 16499 2168 16505 2220
rect 15521 2016 15527 2068
rect 15579 2016 15585 2068
rect 15439 1242 15445 1294
rect 15497 1242 15503 1294
rect 16546 1130 16580 2256
rect 16622 1142 16650 2256
rect 17689 2168 17695 2220
rect 17747 2168 17753 2220
rect 16769 2016 16775 2068
rect 16827 2016 16833 2068
rect 16687 1242 16693 1294
rect 16745 1242 16751 1294
rect 17794 1130 17828 2256
rect 17870 1142 17898 2256
rect 18937 2168 18943 2220
rect 18995 2168 19001 2220
rect 18017 2016 18023 2068
rect 18075 2016 18081 2068
rect 17935 1242 17941 1294
rect 17993 1242 17999 1294
rect 19042 1130 19076 2256
rect 19118 1142 19146 2256
rect 20185 2168 20191 2220
rect 20243 2168 20249 2220
rect 19265 2016 19271 2068
rect 19323 2016 19329 2068
rect 19183 1242 19189 1294
rect 19241 1242 19247 1294
rect 20290 1130 20324 2256
rect 20366 1142 20394 2256
rect 21433 2168 21439 2220
rect 21491 2168 21497 2220
rect 20513 2016 20519 2068
rect 20571 2016 20577 2068
rect 20431 1242 20437 1294
rect 20489 1242 20495 1294
rect 21538 1130 21572 2256
rect 21614 1142 21642 2256
rect 22681 2168 22687 2220
rect 22739 2168 22745 2220
rect 21761 2016 21767 2068
rect 21819 2016 21825 2068
rect 21679 1242 21685 1294
rect 21737 1242 21743 1294
rect 22786 1130 22820 2256
rect 22862 1142 22890 2256
rect 23929 2168 23935 2220
rect 23987 2168 23993 2220
rect 23009 2016 23015 2068
rect 23067 2016 23073 2068
rect 22927 1242 22933 1294
rect 22985 1242 22991 1294
rect 24034 1130 24068 2256
rect 24110 1142 24138 2256
rect 25177 2168 25183 2220
rect 25235 2168 25241 2220
rect 24257 2016 24263 2068
rect 24315 2016 24321 2068
rect 24175 1242 24181 1294
rect 24233 1242 24239 1294
rect 25282 1130 25316 2256
rect 25358 1142 25386 2256
rect 26425 2168 26431 2220
rect 26483 2168 26489 2220
rect 25505 2016 25511 2068
rect 25563 2016 25569 2068
rect 25423 1242 25429 1294
rect 25481 1242 25487 1294
rect 26530 1130 26564 2256
rect 26606 1142 26634 2256
rect 27673 2168 27679 2220
rect 27731 2168 27737 2220
rect 26753 2016 26759 2068
rect 26811 2016 26817 2068
rect 26671 1242 26677 1294
rect 26729 1242 26735 1294
rect 27778 1130 27812 2256
rect 27854 1142 27882 2256
rect 28921 2168 28927 2220
rect 28979 2168 28985 2220
rect 28001 2016 28007 2068
rect 28059 2016 28065 2068
rect 27919 1242 27925 1294
rect 27977 1242 27983 1294
rect 29026 1130 29060 2256
rect 29102 1142 29130 2256
rect 30169 2168 30175 2220
rect 30227 2168 30233 2220
rect 29249 2016 29255 2068
rect 29307 2016 29313 2068
rect 29167 1242 29173 1294
rect 29225 1242 29231 1294
rect 30274 1130 30308 2256
rect 30350 1142 30378 2256
rect 31417 2168 31423 2220
rect 31475 2168 31481 2220
rect 30497 2016 30503 2068
rect 30555 2016 30561 2068
rect 30415 1242 30421 1294
rect 30473 1242 30479 1294
rect 31522 1130 31556 2256
rect 31598 1142 31626 2256
rect 32665 2168 32671 2220
rect 32723 2168 32729 2220
rect 31745 2016 31751 2068
rect 31803 2016 31809 2068
rect 31663 1242 31669 1294
rect 31721 1242 31727 1294
rect 32770 1130 32804 2256
rect 32846 1142 32874 2256
rect 33913 2168 33919 2220
rect 33971 2168 33977 2220
rect 32993 2016 32999 2068
rect 33051 2016 33057 2068
rect 32911 1242 32917 1294
rect 32969 1242 32975 1294
rect 34018 1130 34052 2256
rect 34094 1142 34122 2256
rect 35161 2168 35167 2220
rect 35219 2168 35225 2220
rect 34241 2016 34247 2068
rect 34299 2016 34305 2068
rect 34159 1242 34165 1294
rect 34217 1242 34223 1294
rect 35266 1130 35300 2256
rect 35342 1142 35370 2256
rect 36409 2168 36415 2220
rect 36467 2168 36473 2220
rect 35489 2016 35495 2068
rect 35547 2016 35553 2068
rect 35407 1242 35413 1294
rect 35465 1242 35471 1294
rect 36514 1130 36548 2256
rect 36590 1142 36618 2256
rect 37657 2168 37663 2220
rect 37715 2168 37721 2220
rect 36737 2016 36743 2068
rect 36795 2016 36801 2068
rect 36655 1242 36661 1294
rect 36713 1242 36719 1294
rect 37762 1130 37796 2256
rect 37838 1142 37866 2256
rect 38905 2168 38911 2220
rect 38963 2168 38969 2220
rect 37985 2016 37991 2068
rect 38043 2016 38049 2068
rect 37903 1242 37909 1294
rect 37961 1242 37967 1294
rect 39010 1130 39044 2256
rect 39086 1142 39114 2256
rect 40153 2168 40159 2220
rect 40211 2168 40217 2220
rect 39233 2016 39239 2068
rect 39291 2016 39297 2068
rect 39151 1242 39157 1294
rect 39209 1242 39215 1294
rect 40258 1130 40292 2256
rect 40334 1142 40362 2256
rect 40481 2016 40487 2068
rect 40539 2016 40545 2068
rect 40399 1242 40405 1294
rect 40457 1242 40463 1294
rect 1723 404 1729 456
rect 1781 404 1787 456
rect 2971 404 2977 456
rect 3029 404 3035 456
rect 4219 404 4225 456
rect 4277 404 4283 456
rect 5467 404 5473 456
rect 5525 404 5531 456
rect 6715 404 6721 456
rect 6773 404 6779 456
rect 7963 404 7969 456
rect 8021 404 8027 456
rect 9211 404 9217 456
rect 9269 404 9275 456
rect 10459 404 10465 456
rect 10517 404 10523 456
rect 11707 404 11713 456
rect 11765 404 11771 456
rect 12955 404 12961 456
rect 13013 404 13019 456
rect 14203 404 14209 456
rect 14261 404 14267 456
rect 15451 404 15457 456
rect 15509 404 15515 456
rect 16699 404 16705 456
rect 16757 404 16763 456
rect 17947 404 17953 456
rect 18005 404 18011 456
rect 19195 404 19201 456
rect 19253 404 19259 456
rect 20443 404 20449 456
rect 20501 404 20507 456
rect 21691 404 21697 456
rect 21749 404 21755 456
rect 22939 404 22945 456
rect 22997 404 23003 456
rect 24187 404 24193 456
rect 24245 404 24251 456
rect 25435 404 25441 456
rect 25493 404 25499 456
rect 26683 404 26689 456
rect 26741 404 26747 456
rect 27931 404 27937 456
rect 27989 404 27995 456
rect 29179 404 29185 456
rect 29237 404 29243 456
rect 30427 404 30433 456
rect 30485 404 30491 456
rect 31675 404 31681 456
rect 31733 404 31739 456
rect 32923 404 32929 456
rect 32981 404 32987 456
rect 34171 404 34177 456
rect 34229 404 34235 456
rect 35419 404 35425 456
rect 35477 404 35483 456
rect 36667 404 36673 456
rect 36725 404 36731 456
rect 37915 404 37921 456
rect 37973 404 37979 456
rect 39163 404 39169 456
rect 39221 404 39227 456
rect 40411 404 40417 456
rect 40469 404 40475 456
rect 1478 0 1524 254
rect 1723 82 1729 134
rect 1781 82 1787 134
rect 2726 0 2772 254
rect 2971 82 2977 134
rect 3029 82 3035 134
rect 3974 0 4020 254
rect 4219 82 4225 134
rect 4277 82 4283 134
rect 5222 0 5268 254
rect 5467 82 5473 134
rect 5525 82 5531 134
rect 6470 0 6516 254
rect 6715 82 6721 134
rect 6773 82 6779 134
rect 7718 0 7764 254
rect 7963 82 7969 134
rect 8021 82 8027 134
rect 8966 0 9012 254
rect 9211 82 9217 134
rect 9269 82 9275 134
rect 10214 0 10260 254
rect 10459 82 10465 134
rect 10517 82 10523 134
rect 11462 0 11508 254
rect 11707 82 11713 134
rect 11765 82 11771 134
rect 12710 0 12756 254
rect 12955 82 12961 134
rect 13013 82 13019 134
rect 13958 0 14004 254
rect 14203 82 14209 134
rect 14261 82 14267 134
rect 15206 0 15252 254
rect 15451 82 15457 134
rect 15509 82 15515 134
rect 16454 0 16500 254
rect 16699 82 16705 134
rect 16757 82 16763 134
rect 17702 0 17748 254
rect 17947 82 17953 134
rect 18005 82 18011 134
rect 18950 0 18996 254
rect 19195 82 19201 134
rect 19253 82 19259 134
rect 20198 0 20244 254
rect 20443 82 20449 134
rect 20501 82 20507 134
rect 21446 0 21492 254
rect 21691 82 21697 134
rect 21749 82 21755 134
rect 22694 0 22740 254
rect 22939 82 22945 134
rect 22997 82 23003 134
rect 23942 0 23988 254
rect 24187 82 24193 134
rect 24245 82 24251 134
rect 25190 0 25236 254
rect 25435 82 25441 134
rect 25493 82 25499 134
rect 26438 0 26484 254
rect 26683 82 26689 134
rect 26741 82 26747 134
rect 27686 0 27732 254
rect 27931 82 27937 134
rect 27989 82 27995 134
rect 28934 0 28980 254
rect 29179 82 29185 134
rect 29237 82 29243 134
rect 30182 0 30228 254
rect 30427 82 30433 134
rect 30485 82 30491 134
rect 31430 0 31476 254
rect 31675 82 31681 134
rect 31733 82 31739 134
rect 32678 0 32724 254
rect 32923 82 32929 134
rect 32981 82 32987 134
rect 33926 0 33972 254
rect 34171 82 34177 134
rect 34229 82 34235 134
rect 35174 0 35220 254
rect 35419 82 35425 134
rect 35477 82 35483 134
rect 36422 0 36468 254
rect 36667 82 36673 134
rect 36725 82 36731 134
rect 37670 0 37716 254
rect 37915 82 37921 134
rect 37973 82 37979 134
rect 38918 0 38964 254
rect 39163 82 39169 134
rect 39221 82 39227 134
rect 40166 0 40212 254
rect 40411 82 40417 134
rect 40469 82 40475 134
<< via1 >>
rect 1471 2168 1523 2220
rect 2719 2168 2771 2220
rect 1799 2016 1851 2068
rect 1717 1242 1769 1294
rect 3967 2168 4019 2220
rect 3047 2016 3099 2068
rect 2965 1242 3017 1294
rect 5215 2168 5267 2220
rect 4295 2016 4347 2068
rect 4213 1242 4265 1294
rect 6463 2168 6515 2220
rect 5543 2016 5595 2068
rect 5461 1242 5513 1294
rect 7711 2168 7763 2220
rect 6791 2016 6843 2068
rect 6709 1242 6761 1294
rect 8959 2168 9011 2220
rect 8039 2016 8091 2068
rect 7957 1242 8009 1294
rect 10207 2168 10259 2220
rect 9287 2016 9339 2068
rect 9205 1242 9257 1294
rect 11455 2168 11507 2220
rect 10535 2016 10587 2068
rect 10453 1242 10505 1294
rect 12703 2168 12755 2220
rect 11783 2016 11835 2068
rect 11701 1242 11753 1294
rect 13951 2168 14003 2220
rect 13031 2016 13083 2068
rect 12949 1242 13001 1294
rect 15199 2168 15251 2220
rect 14279 2016 14331 2068
rect 14197 1242 14249 1294
rect 16447 2168 16499 2220
rect 15527 2016 15579 2068
rect 15445 1242 15497 1294
rect 17695 2168 17747 2220
rect 16775 2016 16827 2068
rect 16693 1242 16745 1294
rect 18943 2168 18995 2220
rect 18023 2016 18075 2068
rect 17941 1242 17993 1294
rect 20191 2168 20243 2220
rect 19271 2016 19323 2068
rect 19189 1242 19241 1294
rect 21439 2168 21491 2220
rect 20519 2016 20571 2068
rect 20437 1242 20489 1294
rect 22687 2168 22739 2220
rect 21767 2016 21819 2068
rect 21685 1242 21737 1294
rect 23935 2168 23987 2220
rect 23015 2016 23067 2068
rect 22933 1242 22985 1294
rect 25183 2168 25235 2220
rect 24263 2016 24315 2068
rect 24181 1242 24233 1294
rect 26431 2168 26483 2220
rect 25511 2016 25563 2068
rect 25429 1242 25481 1294
rect 27679 2168 27731 2220
rect 26759 2016 26811 2068
rect 26677 1242 26729 1294
rect 28927 2168 28979 2220
rect 28007 2016 28059 2068
rect 27925 1242 27977 1294
rect 30175 2168 30227 2220
rect 29255 2016 29307 2068
rect 29173 1242 29225 1294
rect 31423 2168 31475 2220
rect 30503 2016 30555 2068
rect 30421 1242 30473 1294
rect 32671 2168 32723 2220
rect 31751 2016 31803 2068
rect 31669 1242 31721 1294
rect 33919 2168 33971 2220
rect 32999 2016 33051 2068
rect 32917 1242 32969 1294
rect 35167 2168 35219 2220
rect 34247 2016 34299 2068
rect 34165 1242 34217 1294
rect 36415 2168 36467 2220
rect 35495 2016 35547 2068
rect 35413 1242 35465 1294
rect 37663 2168 37715 2220
rect 36743 2016 36795 2068
rect 36661 1242 36713 1294
rect 38911 2168 38963 2220
rect 37991 2016 38043 2068
rect 37909 1242 37961 1294
rect 40159 2168 40211 2220
rect 39239 2016 39291 2068
rect 39157 1242 39209 1294
rect 40487 2016 40539 2068
rect 40405 1242 40457 1294
rect 1729 404 1781 456
rect 2977 404 3029 456
rect 4225 404 4277 456
rect 5473 404 5525 456
rect 6721 404 6773 456
rect 7969 404 8021 456
rect 9217 404 9269 456
rect 10465 404 10517 456
rect 11713 404 11765 456
rect 12961 404 13013 456
rect 14209 404 14261 456
rect 15457 404 15509 456
rect 16705 404 16757 456
rect 17953 404 18005 456
rect 19201 404 19253 456
rect 20449 404 20501 456
rect 21697 404 21749 456
rect 22945 404 22997 456
rect 24193 404 24245 456
rect 25441 404 25493 456
rect 26689 404 26741 456
rect 27937 404 27989 456
rect 29185 404 29237 456
rect 30433 404 30485 456
rect 31681 404 31733 456
rect 32929 404 32981 456
rect 34177 404 34229 456
rect 35425 404 35477 456
rect 36673 404 36725 456
rect 37921 404 37973 456
rect 39169 404 39221 456
rect 40417 404 40469 456
rect 1729 82 1781 134
rect 2977 82 3029 134
rect 4225 82 4277 134
rect 5473 82 5525 134
rect 6721 82 6773 134
rect 7969 82 8021 134
rect 9217 82 9269 134
rect 10465 82 10517 134
rect 11713 82 11765 134
rect 12961 82 13013 134
rect 14209 82 14261 134
rect 15457 82 15509 134
rect 16705 82 16757 134
rect 17953 82 18005 134
rect 19201 82 19253 134
rect 20449 82 20501 134
rect 21697 82 21749 134
rect 22945 82 22997 134
rect 24193 82 24245 134
rect 25441 82 25493 134
rect 26689 82 26741 134
rect 27937 82 27989 134
rect 29185 82 29237 134
rect 30433 82 30485 134
rect 31681 82 31733 134
rect 32929 82 32981 134
rect 34177 82 34229 134
rect 35425 82 35477 134
rect 36673 82 36725 134
rect 37921 82 37973 134
rect 39169 82 39221 134
rect 40417 82 40469 134
<< metal2 >>
rect 1469 2222 1525 2231
rect 1469 2157 1525 2166
rect 2717 2222 2773 2231
rect 2717 2157 2773 2166
rect 3965 2222 4021 2231
rect 3965 2157 4021 2166
rect 5213 2222 5269 2231
rect 5213 2157 5269 2166
rect 6461 2222 6517 2231
rect 6461 2157 6517 2166
rect 7709 2222 7765 2231
rect 7709 2157 7765 2166
rect 8957 2222 9013 2231
rect 8957 2157 9013 2166
rect 10205 2222 10261 2231
rect 10205 2157 10261 2166
rect 11453 2222 11509 2231
rect 11453 2157 11509 2166
rect 12701 2222 12757 2231
rect 12701 2157 12757 2166
rect 13949 2222 14005 2231
rect 13949 2157 14005 2166
rect 15197 2222 15253 2231
rect 15197 2157 15253 2166
rect 16445 2222 16501 2231
rect 16445 2157 16501 2166
rect 17693 2222 17749 2231
rect 17693 2157 17749 2166
rect 18941 2222 18997 2231
rect 18941 2157 18997 2166
rect 20189 2222 20245 2231
rect 20189 2157 20245 2166
rect 21437 2222 21493 2231
rect 21437 2157 21493 2166
rect 22685 2222 22741 2231
rect 22685 2157 22741 2166
rect 23933 2222 23989 2231
rect 23933 2157 23989 2166
rect 25181 2222 25237 2231
rect 25181 2157 25237 2166
rect 26429 2222 26485 2231
rect 26429 2157 26485 2166
rect 27677 2222 27733 2231
rect 27677 2157 27733 2166
rect 28925 2222 28981 2231
rect 28925 2157 28981 2166
rect 30173 2222 30229 2231
rect 30173 2157 30229 2166
rect 31421 2222 31477 2231
rect 31421 2157 31477 2166
rect 32669 2222 32725 2231
rect 32669 2157 32725 2166
rect 33917 2222 33973 2231
rect 33917 2157 33973 2166
rect 35165 2222 35221 2231
rect 35165 2157 35221 2166
rect 36413 2222 36469 2231
rect 36413 2157 36469 2166
rect 37661 2222 37717 2231
rect 37661 2157 37717 2166
rect 38909 2222 38965 2231
rect 38909 2157 38965 2166
rect 40157 2222 40213 2231
rect 40157 2157 40213 2166
rect 1797 2070 1853 2079
rect 1797 2005 1853 2014
rect 3045 2070 3101 2079
rect 3045 2005 3101 2014
rect 4293 2070 4349 2079
rect 4293 2005 4349 2014
rect 5541 2070 5597 2079
rect 5541 2005 5597 2014
rect 6789 2070 6845 2079
rect 6789 2005 6845 2014
rect 8037 2070 8093 2079
rect 8037 2005 8093 2014
rect 9285 2070 9341 2079
rect 9285 2005 9341 2014
rect 10533 2070 10589 2079
rect 10533 2005 10589 2014
rect 11781 2070 11837 2079
rect 11781 2005 11837 2014
rect 13029 2070 13085 2079
rect 13029 2005 13085 2014
rect 14277 2070 14333 2079
rect 14277 2005 14333 2014
rect 15525 2070 15581 2079
rect 15525 2005 15581 2014
rect 16773 2070 16829 2079
rect 16773 2005 16829 2014
rect 18021 2070 18077 2079
rect 18021 2005 18077 2014
rect 19269 2070 19325 2079
rect 19269 2005 19325 2014
rect 20517 2070 20573 2079
rect 20517 2005 20573 2014
rect 21765 2070 21821 2079
rect 21765 2005 21821 2014
rect 23013 2070 23069 2079
rect 23013 2005 23069 2014
rect 24261 2070 24317 2079
rect 24261 2005 24317 2014
rect 25509 2070 25565 2079
rect 25509 2005 25565 2014
rect 26757 2070 26813 2079
rect 26757 2005 26813 2014
rect 28005 2070 28061 2079
rect 28005 2005 28061 2014
rect 29253 2070 29309 2079
rect 29253 2005 29309 2014
rect 30501 2070 30557 2079
rect 30501 2005 30557 2014
rect 31749 2070 31805 2079
rect 31749 2005 31805 2014
rect 32997 2070 33053 2079
rect 32997 2005 33053 2014
rect 34245 2070 34301 2079
rect 34245 2005 34301 2014
rect 35493 2070 35549 2079
rect 35493 2005 35549 2014
rect 36741 2070 36797 2079
rect 36741 2005 36797 2014
rect 37989 2070 38045 2079
rect 37989 2005 38045 2014
rect 39237 2070 39293 2079
rect 39237 2005 39293 2014
rect 40485 2070 40541 2079
rect 40485 2005 40541 2014
rect 1715 1296 1771 1305
rect 1715 1231 1771 1240
rect 2963 1296 3019 1305
rect 2963 1231 3019 1240
rect 4211 1296 4267 1305
rect 4211 1231 4267 1240
rect 5459 1296 5515 1305
rect 5459 1231 5515 1240
rect 6707 1296 6763 1305
rect 6707 1231 6763 1240
rect 7955 1296 8011 1305
rect 7955 1231 8011 1240
rect 9203 1296 9259 1305
rect 9203 1231 9259 1240
rect 10451 1296 10507 1305
rect 10451 1231 10507 1240
rect 11699 1296 11755 1305
rect 11699 1231 11755 1240
rect 12947 1296 13003 1305
rect 12947 1231 13003 1240
rect 14195 1296 14251 1305
rect 14195 1231 14251 1240
rect 15443 1296 15499 1305
rect 15443 1231 15499 1240
rect 16691 1296 16747 1305
rect 16691 1231 16747 1240
rect 17939 1296 17995 1305
rect 17939 1231 17995 1240
rect 19187 1296 19243 1305
rect 19187 1231 19243 1240
rect 20435 1296 20491 1305
rect 20435 1231 20491 1240
rect 21683 1296 21739 1305
rect 21683 1231 21739 1240
rect 22931 1296 22987 1305
rect 22931 1231 22987 1240
rect 24179 1296 24235 1305
rect 24179 1231 24235 1240
rect 25427 1296 25483 1305
rect 25427 1231 25483 1240
rect 26675 1296 26731 1305
rect 26675 1231 26731 1240
rect 27923 1296 27979 1305
rect 27923 1231 27979 1240
rect 29171 1296 29227 1305
rect 29171 1231 29227 1240
rect 30419 1296 30475 1305
rect 30419 1231 30475 1240
rect 31667 1296 31723 1305
rect 31667 1231 31723 1240
rect 32915 1296 32971 1305
rect 32915 1231 32971 1240
rect 34163 1296 34219 1305
rect 34163 1231 34219 1240
rect 35411 1296 35467 1305
rect 35411 1231 35467 1240
rect 36659 1296 36715 1305
rect 36659 1231 36715 1240
rect 37907 1296 37963 1305
rect 37907 1231 37963 1240
rect 39155 1296 39211 1305
rect 39155 1231 39211 1240
rect 40403 1296 40459 1305
rect 40403 1231 40459 1240
rect 1727 458 1783 467
rect 1727 393 1783 402
rect 2975 458 3031 467
rect 2975 393 3031 402
rect 4223 458 4279 467
rect 4223 393 4279 402
rect 5471 458 5527 467
rect 5471 393 5527 402
rect 6719 458 6775 467
rect 6719 393 6775 402
rect 7967 458 8023 467
rect 7967 393 8023 402
rect 9215 458 9271 467
rect 9215 393 9271 402
rect 10463 458 10519 467
rect 10463 393 10519 402
rect 11711 458 11767 467
rect 11711 393 11767 402
rect 12959 458 13015 467
rect 12959 393 13015 402
rect 14207 458 14263 467
rect 14207 393 14263 402
rect 15455 458 15511 467
rect 15455 393 15511 402
rect 16703 458 16759 467
rect 16703 393 16759 402
rect 17951 458 18007 467
rect 17951 393 18007 402
rect 19199 458 19255 467
rect 19199 393 19255 402
rect 20447 458 20503 467
rect 20447 393 20503 402
rect 21695 458 21751 467
rect 21695 393 21751 402
rect 22943 458 22999 467
rect 22943 393 22999 402
rect 24191 458 24247 467
rect 24191 393 24247 402
rect 25439 458 25495 467
rect 25439 393 25495 402
rect 26687 458 26743 467
rect 26687 393 26743 402
rect 27935 458 27991 467
rect 27935 393 27991 402
rect 29183 458 29239 467
rect 29183 393 29239 402
rect 30431 458 30487 467
rect 30431 393 30487 402
rect 31679 458 31735 467
rect 31679 393 31735 402
rect 32927 458 32983 467
rect 32927 393 32983 402
rect 34175 458 34231 467
rect 34175 393 34231 402
rect 35423 458 35479 467
rect 35423 393 35479 402
rect 36671 458 36727 467
rect 36671 393 36727 402
rect 37919 458 37975 467
rect 37919 393 37975 402
rect 39167 458 39223 467
rect 39167 393 39223 402
rect 40415 458 40471 467
rect 40415 393 40471 402
rect 1727 136 1783 145
rect 1727 71 1783 80
rect 2975 136 3031 145
rect 2975 71 3031 80
rect 4223 136 4279 145
rect 4223 71 4279 80
rect 5471 136 5527 145
rect 5471 71 5527 80
rect 6719 136 6775 145
rect 6719 71 6775 80
rect 7967 136 8023 145
rect 7967 71 8023 80
rect 9215 136 9271 145
rect 9215 71 9271 80
rect 10463 136 10519 145
rect 10463 71 10519 80
rect 11711 136 11767 145
rect 11711 71 11767 80
rect 12959 136 13015 145
rect 12959 71 13015 80
rect 14207 136 14263 145
rect 14207 71 14263 80
rect 15455 136 15511 145
rect 15455 71 15511 80
rect 16703 136 16759 145
rect 16703 71 16759 80
rect 17951 136 18007 145
rect 17951 71 18007 80
rect 19199 136 19255 145
rect 19199 71 19255 80
rect 20447 136 20503 145
rect 20447 71 20503 80
rect 21695 136 21751 145
rect 21695 71 21751 80
rect 22943 136 22999 145
rect 22943 71 22999 80
rect 24191 136 24247 145
rect 24191 71 24247 80
rect 25439 136 25495 145
rect 25439 71 25495 80
rect 26687 136 26743 145
rect 26687 71 26743 80
rect 27935 136 27991 145
rect 27935 71 27991 80
rect 29183 136 29239 145
rect 29183 71 29239 80
rect 30431 136 30487 145
rect 30431 71 30487 80
rect 31679 136 31735 145
rect 31679 71 31735 80
rect 32927 136 32983 145
rect 32927 71 32983 80
rect 34175 136 34231 145
rect 34175 71 34231 80
rect 35423 136 35479 145
rect 35423 71 35479 80
rect 36671 136 36727 145
rect 36671 71 36727 80
rect 37919 136 37975 145
rect 37919 71 37975 80
rect 39167 136 39223 145
rect 39167 71 39223 80
rect 40415 136 40471 145
rect 40415 71 40471 80
<< via2 >>
rect 1469 2220 1525 2222
rect 1469 2168 1471 2220
rect 1471 2168 1523 2220
rect 1523 2168 1525 2220
rect 1469 2166 1525 2168
rect 2717 2220 2773 2222
rect 2717 2168 2719 2220
rect 2719 2168 2771 2220
rect 2771 2168 2773 2220
rect 2717 2166 2773 2168
rect 3965 2220 4021 2222
rect 3965 2168 3967 2220
rect 3967 2168 4019 2220
rect 4019 2168 4021 2220
rect 3965 2166 4021 2168
rect 5213 2220 5269 2222
rect 5213 2168 5215 2220
rect 5215 2168 5267 2220
rect 5267 2168 5269 2220
rect 5213 2166 5269 2168
rect 6461 2220 6517 2222
rect 6461 2168 6463 2220
rect 6463 2168 6515 2220
rect 6515 2168 6517 2220
rect 6461 2166 6517 2168
rect 7709 2220 7765 2222
rect 7709 2168 7711 2220
rect 7711 2168 7763 2220
rect 7763 2168 7765 2220
rect 7709 2166 7765 2168
rect 8957 2220 9013 2222
rect 8957 2168 8959 2220
rect 8959 2168 9011 2220
rect 9011 2168 9013 2220
rect 8957 2166 9013 2168
rect 10205 2220 10261 2222
rect 10205 2168 10207 2220
rect 10207 2168 10259 2220
rect 10259 2168 10261 2220
rect 10205 2166 10261 2168
rect 11453 2220 11509 2222
rect 11453 2168 11455 2220
rect 11455 2168 11507 2220
rect 11507 2168 11509 2220
rect 11453 2166 11509 2168
rect 12701 2220 12757 2222
rect 12701 2168 12703 2220
rect 12703 2168 12755 2220
rect 12755 2168 12757 2220
rect 12701 2166 12757 2168
rect 13949 2220 14005 2222
rect 13949 2168 13951 2220
rect 13951 2168 14003 2220
rect 14003 2168 14005 2220
rect 13949 2166 14005 2168
rect 15197 2220 15253 2222
rect 15197 2168 15199 2220
rect 15199 2168 15251 2220
rect 15251 2168 15253 2220
rect 15197 2166 15253 2168
rect 16445 2220 16501 2222
rect 16445 2168 16447 2220
rect 16447 2168 16499 2220
rect 16499 2168 16501 2220
rect 16445 2166 16501 2168
rect 17693 2220 17749 2222
rect 17693 2168 17695 2220
rect 17695 2168 17747 2220
rect 17747 2168 17749 2220
rect 17693 2166 17749 2168
rect 18941 2220 18997 2222
rect 18941 2168 18943 2220
rect 18943 2168 18995 2220
rect 18995 2168 18997 2220
rect 18941 2166 18997 2168
rect 20189 2220 20245 2222
rect 20189 2168 20191 2220
rect 20191 2168 20243 2220
rect 20243 2168 20245 2220
rect 20189 2166 20245 2168
rect 21437 2220 21493 2222
rect 21437 2168 21439 2220
rect 21439 2168 21491 2220
rect 21491 2168 21493 2220
rect 21437 2166 21493 2168
rect 22685 2220 22741 2222
rect 22685 2168 22687 2220
rect 22687 2168 22739 2220
rect 22739 2168 22741 2220
rect 22685 2166 22741 2168
rect 23933 2220 23989 2222
rect 23933 2168 23935 2220
rect 23935 2168 23987 2220
rect 23987 2168 23989 2220
rect 23933 2166 23989 2168
rect 25181 2220 25237 2222
rect 25181 2168 25183 2220
rect 25183 2168 25235 2220
rect 25235 2168 25237 2220
rect 25181 2166 25237 2168
rect 26429 2220 26485 2222
rect 26429 2168 26431 2220
rect 26431 2168 26483 2220
rect 26483 2168 26485 2220
rect 26429 2166 26485 2168
rect 27677 2220 27733 2222
rect 27677 2168 27679 2220
rect 27679 2168 27731 2220
rect 27731 2168 27733 2220
rect 27677 2166 27733 2168
rect 28925 2220 28981 2222
rect 28925 2168 28927 2220
rect 28927 2168 28979 2220
rect 28979 2168 28981 2220
rect 28925 2166 28981 2168
rect 30173 2220 30229 2222
rect 30173 2168 30175 2220
rect 30175 2168 30227 2220
rect 30227 2168 30229 2220
rect 30173 2166 30229 2168
rect 31421 2220 31477 2222
rect 31421 2168 31423 2220
rect 31423 2168 31475 2220
rect 31475 2168 31477 2220
rect 31421 2166 31477 2168
rect 32669 2220 32725 2222
rect 32669 2168 32671 2220
rect 32671 2168 32723 2220
rect 32723 2168 32725 2220
rect 32669 2166 32725 2168
rect 33917 2220 33973 2222
rect 33917 2168 33919 2220
rect 33919 2168 33971 2220
rect 33971 2168 33973 2220
rect 33917 2166 33973 2168
rect 35165 2220 35221 2222
rect 35165 2168 35167 2220
rect 35167 2168 35219 2220
rect 35219 2168 35221 2220
rect 35165 2166 35221 2168
rect 36413 2220 36469 2222
rect 36413 2168 36415 2220
rect 36415 2168 36467 2220
rect 36467 2168 36469 2220
rect 36413 2166 36469 2168
rect 37661 2220 37717 2222
rect 37661 2168 37663 2220
rect 37663 2168 37715 2220
rect 37715 2168 37717 2220
rect 37661 2166 37717 2168
rect 38909 2220 38965 2222
rect 38909 2168 38911 2220
rect 38911 2168 38963 2220
rect 38963 2168 38965 2220
rect 38909 2166 38965 2168
rect 40157 2220 40213 2222
rect 40157 2168 40159 2220
rect 40159 2168 40211 2220
rect 40211 2168 40213 2220
rect 40157 2166 40213 2168
rect 1797 2068 1853 2070
rect 1797 2016 1799 2068
rect 1799 2016 1851 2068
rect 1851 2016 1853 2068
rect 1797 2014 1853 2016
rect 3045 2068 3101 2070
rect 3045 2016 3047 2068
rect 3047 2016 3099 2068
rect 3099 2016 3101 2068
rect 3045 2014 3101 2016
rect 4293 2068 4349 2070
rect 4293 2016 4295 2068
rect 4295 2016 4347 2068
rect 4347 2016 4349 2068
rect 4293 2014 4349 2016
rect 5541 2068 5597 2070
rect 5541 2016 5543 2068
rect 5543 2016 5595 2068
rect 5595 2016 5597 2068
rect 5541 2014 5597 2016
rect 6789 2068 6845 2070
rect 6789 2016 6791 2068
rect 6791 2016 6843 2068
rect 6843 2016 6845 2068
rect 6789 2014 6845 2016
rect 8037 2068 8093 2070
rect 8037 2016 8039 2068
rect 8039 2016 8091 2068
rect 8091 2016 8093 2068
rect 8037 2014 8093 2016
rect 9285 2068 9341 2070
rect 9285 2016 9287 2068
rect 9287 2016 9339 2068
rect 9339 2016 9341 2068
rect 9285 2014 9341 2016
rect 10533 2068 10589 2070
rect 10533 2016 10535 2068
rect 10535 2016 10587 2068
rect 10587 2016 10589 2068
rect 10533 2014 10589 2016
rect 11781 2068 11837 2070
rect 11781 2016 11783 2068
rect 11783 2016 11835 2068
rect 11835 2016 11837 2068
rect 11781 2014 11837 2016
rect 13029 2068 13085 2070
rect 13029 2016 13031 2068
rect 13031 2016 13083 2068
rect 13083 2016 13085 2068
rect 13029 2014 13085 2016
rect 14277 2068 14333 2070
rect 14277 2016 14279 2068
rect 14279 2016 14331 2068
rect 14331 2016 14333 2068
rect 14277 2014 14333 2016
rect 15525 2068 15581 2070
rect 15525 2016 15527 2068
rect 15527 2016 15579 2068
rect 15579 2016 15581 2068
rect 15525 2014 15581 2016
rect 16773 2068 16829 2070
rect 16773 2016 16775 2068
rect 16775 2016 16827 2068
rect 16827 2016 16829 2068
rect 16773 2014 16829 2016
rect 18021 2068 18077 2070
rect 18021 2016 18023 2068
rect 18023 2016 18075 2068
rect 18075 2016 18077 2068
rect 18021 2014 18077 2016
rect 19269 2068 19325 2070
rect 19269 2016 19271 2068
rect 19271 2016 19323 2068
rect 19323 2016 19325 2068
rect 19269 2014 19325 2016
rect 20517 2068 20573 2070
rect 20517 2016 20519 2068
rect 20519 2016 20571 2068
rect 20571 2016 20573 2068
rect 20517 2014 20573 2016
rect 21765 2068 21821 2070
rect 21765 2016 21767 2068
rect 21767 2016 21819 2068
rect 21819 2016 21821 2068
rect 21765 2014 21821 2016
rect 23013 2068 23069 2070
rect 23013 2016 23015 2068
rect 23015 2016 23067 2068
rect 23067 2016 23069 2068
rect 23013 2014 23069 2016
rect 24261 2068 24317 2070
rect 24261 2016 24263 2068
rect 24263 2016 24315 2068
rect 24315 2016 24317 2068
rect 24261 2014 24317 2016
rect 25509 2068 25565 2070
rect 25509 2016 25511 2068
rect 25511 2016 25563 2068
rect 25563 2016 25565 2068
rect 25509 2014 25565 2016
rect 26757 2068 26813 2070
rect 26757 2016 26759 2068
rect 26759 2016 26811 2068
rect 26811 2016 26813 2068
rect 26757 2014 26813 2016
rect 28005 2068 28061 2070
rect 28005 2016 28007 2068
rect 28007 2016 28059 2068
rect 28059 2016 28061 2068
rect 28005 2014 28061 2016
rect 29253 2068 29309 2070
rect 29253 2016 29255 2068
rect 29255 2016 29307 2068
rect 29307 2016 29309 2068
rect 29253 2014 29309 2016
rect 30501 2068 30557 2070
rect 30501 2016 30503 2068
rect 30503 2016 30555 2068
rect 30555 2016 30557 2068
rect 30501 2014 30557 2016
rect 31749 2068 31805 2070
rect 31749 2016 31751 2068
rect 31751 2016 31803 2068
rect 31803 2016 31805 2068
rect 31749 2014 31805 2016
rect 32997 2068 33053 2070
rect 32997 2016 32999 2068
rect 32999 2016 33051 2068
rect 33051 2016 33053 2068
rect 32997 2014 33053 2016
rect 34245 2068 34301 2070
rect 34245 2016 34247 2068
rect 34247 2016 34299 2068
rect 34299 2016 34301 2068
rect 34245 2014 34301 2016
rect 35493 2068 35549 2070
rect 35493 2016 35495 2068
rect 35495 2016 35547 2068
rect 35547 2016 35549 2068
rect 35493 2014 35549 2016
rect 36741 2068 36797 2070
rect 36741 2016 36743 2068
rect 36743 2016 36795 2068
rect 36795 2016 36797 2068
rect 36741 2014 36797 2016
rect 37989 2068 38045 2070
rect 37989 2016 37991 2068
rect 37991 2016 38043 2068
rect 38043 2016 38045 2068
rect 37989 2014 38045 2016
rect 39237 2068 39293 2070
rect 39237 2016 39239 2068
rect 39239 2016 39291 2068
rect 39291 2016 39293 2068
rect 39237 2014 39293 2016
rect 40485 2068 40541 2070
rect 40485 2016 40487 2068
rect 40487 2016 40539 2068
rect 40539 2016 40541 2068
rect 40485 2014 40541 2016
rect 1715 1294 1771 1296
rect 1715 1242 1717 1294
rect 1717 1242 1769 1294
rect 1769 1242 1771 1294
rect 1715 1240 1771 1242
rect 2963 1294 3019 1296
rect 2963 1242 2965 1294
rect 2965 1242 3017 1294
rect 3017 1242 3019 1294
rect 2963 1240 3019 1242
rect 4211 1294 4267 1296
rect 4211 1242 4213 1294
rect 4213 1242 4265 1294
rect 4265 1242 4267 1294
rect 4211 1240 4267 1242
rect 5459 1294 5515 1296
rect 5459 1242 5461 1294
rect 5461 1242 5513 1294
rect 5513 1242 5515 1294
rect 5459 1240 5515 1242
rect 6707 1294 6763 1296
rect 6707 1242 6709 1294
rect 6709 1242 6761 1294
rect 6761 1242 6763 1294
rect 6707 1240 6763 1242
rect 7955 1294 8011 1296
rect 7955 1242 7957 1294
rect 7957 1242 8009 1294
rect 8009 1242 8011 1294
rect 7955 1240 8011 1242
rect 9203 1294 9259 1296
rect 9203 1242 9205 1294
rect 9205 1242 9257 1294
rect 9257 1242 9259 1294
rect 9203 1240 9259 1242
rect 10451 1294 10507 1296
rect 10451 1242 10453 1294
rect 10453 1242 10505 1294
rect 10505 1242 10507 1294
rect 10451 1240 10507 1242
rect 11699 1294 11755 1296
rect 11699 1242 11701 1294
rect 11701 1242 11753 1294
rect 11753 1242 11755 1294
rect 11699 1240 11755 1242
rect 12947 1294 13003 1296
rect 12947 1242 12949 1294
rect 12949 1242 13001 1294
rect 13001 1242 13003 1294
rect 12947 1240 13003 1242
rect 14195 1294 14251 1296
rect 14195 1242 14197 1294
rect 14197 1242 14249 1294
rect 14249 1242 14251 1294
rect 14195 1240 14251 1242
rect 15443 1294 15499 1296
rect 15443 1242 15445 1294
rect 15445 1242 15497 1294
rect 15497 1242 15499 1294
rect 15443 1240 15499 1242
rect 16691 1294 16747 1296
rect 16691 1242 16693 1294
rect 16693 1242 16745 1294
rect 16745 1242 16747 1294
rect 16691 1240 16747 1242
rect 17939 1294 17995 1296
rect 17939 1242 17941 1294
rect 17941 1242 17993 1294
rect 17993 1242 17995 1294
rect 17939 1240 17995 1242
rect 19187 1294 19243 1296
rect 19187 1242 19189 1294
rect 19189 1242 19241 1294
rect 19241 1242 19243 1294
rect 19187 1240 19243 1242
rect 20435 1294 20491 1296
rect 20435 1242 20437 1294
rect 20437 1242 20489 1294
rect 20489 1242 20491 1294
rect 20435 1240 20491 1242
rect 21683 1294 21739 1296
rect 21683 1242 21685 1294
rect 21685 1242 21737 1294
rect 21737 1242 21739 1294
rect 21683 1240 21739 1242
rect 22931 1294 22987 1296
rect 22931 1242 22933 1294
rect 22933 1242 22985 1294
rect 22985 1242 22987 1294
rect 22931 1240 22987 1242
rect 24179 1294 24235 1296
rect 24179 1242 24181 1294
rect 24181 1242 24233 1294
rect 24233 1242 24235 1294
rect 24179 1240 24235 1242
rect 25427 1294 25483 1296
rect 25427 1242 25429 1294
rect 25429 1242 25481 1294
rect 25481 1242 25483 1294
rect 25427 1240 25483 1242
rect 26675 1294 26731 1296
rect 26675 1242 26677 1294
rect 26677 1242 26729 1294
rect 26729 1242 26731 1294
rect 26675 1240 26731 1242
rect 27923 1294 27979 1296
rect 27923 1242 27925 1294
rect 27925 1242 27977 1294
rect 27977 1242 27979 1294
rect 27923 1240 27979 1242
rect 29171 1294 29227 1296
rect 29171 1242 29173 1294
rect 29173 1242 29225 1294
rect 29225 1242 29227 1294
rect 29171 1240 29227 1242
rect 30419 1294 30475 1296
rect 30419 1242 30421 1294
rect 30421 1242 30473 1294
rect 30473 1242 30475 1294
rect 30419 1240 30475 1242
rect 31667 1294 31723 1296
rect 31667 1242 31669 1294
rect 31669 1242 31721 1294
rect 31721 1242 31723 1294
rect 31667 1240 31723 1242
rect 32915 1294 32971 1296
rect 32915 1242 32917 1294
rect 32917 1242 32969 1294
rect 32969 1242 32971 1294
rect 32915 1240 32971 1242
rect 34163 1294 34219 1296
rect 34163 1242 34165 1294
rect 34165 1242 34217 1294
rect 34217 1242 34219 1294
rect 34163 1240 34219 1242
rect 35411 1294 35467 1296
rect 35411 1242 35413 1294
rect 35413 1242 35465 1294
rect 35465 1242 35467 1294
rect 35411 1240 35467 1242
rect 36659 1294 36715 1296
rect 36659 1242 36661 1294
rect 36661 1242 36713 1294
rect 36713 1242 36715 1294
rect 36659 1240 36715 1242
rect 37907 1294 37963 1296
rect 37907 1242 37909 1294
rect 37909 1242 37961 1294
rect 37961 1242 37963 1294
rect 37907 1240 37963 1242
rect 39155 1294 39211 1296
rect 39155 1242 39157 1294
rect 39157 1242 39209 1294
rect 39209 1242 39211 1294
rect 39155 1240 39211 1242
rect 40403 1294 40459 1296
rect 40403 1242 40405 1294
rect 40405 1242 40457 1294
rect 40457 1242 40459 1294
rect 40403 1240 40459 1242
rect 1727 456 1783 458
rect 1727 404 1729 456
rect 1729 404 1781 456
rect 1781 404 1783 456
rect 1727 402 1783 404
rect 2975 456 3031 458
rect 2975 404 2977 456
rect 2977 404 3029 456
rect 3029 404 3031 456
rect 2975 402 3031 404
rect 4223 456 4279 458
rect 4223 404 4225 456
rect 4225 404 4277 456
rect 4277 404 4279 456
rect 4223 402 4279 404
rect 5471 456 5527 458
rect 5471 404 5473 456
rect 5473 404 5525 456
rect 5525 404 5527 456
rect 5471 402 5527 404
rect 6719 456 6775 458
rect 6719 404 6721 456
rect 6721 404 6773 456
rect 6773 404 6775 456
rect 6719 402 6775 404
rect 7967 456 8023 458
rect 7967 404 7969 456
rect 7969 404 8021 456
rect 8021 404 8023 456
rect 7967 402 8023 404
rect 9215 456 9271 458
rect 9215 404 9217 456
rect 9217 404 9269 456
rect 9269 404 9271 456
rect 9215 402 9271 404
rect 10463 456 10519 458
rect 10463 404 10465 456
rect 10465 404 10517 456
rect 10517 404 10519 456
rect 10463 402 10519 404
rect 11711 456 11767 458
rect 11711 404 11713 456
rect 11713 404 11765 456
rect 11765 404 11767 456
rect 11711 402 11767 404
rect 12959 456 13015 458
rect 12959 404 12961 456
rect 12961 404 13013 456
rect 13013 404 13015 456
rect 12959 402 13015 404
rect 14207 456 14263 458
rect 14207 404 14209 456
rect 14209 404 14261 456
rect 14261 404 14263 456
rect 14207 402 14263 404
rect 15455 456 15511 458
rect 15455 404 15457 456
rect 15457 404 15509 456
rect 15509 404 15511 456
rect 15455 402 15511 404
rect 16703 456 16759 458
rect 16703 404 16705 456
rect 16705 404 16757 456
rect 16757 404 16759 456
rect 16703 402 16759 404
rect 17951 456 18007 458
rect 17951 404 17953 456
rect 17953 404 18005 456
rect 18005 404 18007 456
rect 17951 402 18007 404
rect 19199 456 19255 458
rect 19199 404 19201 456
rect 19201 404 19253 456
rect 19253 404 19255 456
rect 19199 402 19255 404
rect 20447 456 20503 458
rect 20447 404 20449 456
rect 20449 404 20501 456
rect 20501 404 20503 456
rect 20447 402 20503 404
rect 21695 456 21751 458
rect 21695 404 21697 456
rect 21697 404 21749 456
rect 21749 404 21751 456
rect 21695 402 21751 404
rect 22943 456 22999 458
rect 22943 404 22945 456
rect 22945 404 22997 456
rect 22997 404 22999 456
rect 22943 402 22999 404
rect 24191 456 24247 458
rect 24191 404 24193 456
rect 24193 404 24245 456
rect 24245 404 24247 456
rect 24191 402 24247 404
rect 25439 456 25495 458
rect 25439 404 25441 456
rect 25441 404 25493 456
rect 25493 404 25495 456
rect 25439 402 25495 404
rect 26687 456 26743 458
rect 26687 404 26689 456
rect 26689 404 26741 456
rect 26741 404 26743 456
rect 26687 402 26743 404
rect 27935 456 27991 458
rect 27935 404 27937 456
rect 27937 404 27989 456
rect 27989 404 27991 456
rect 27935 402 27991 404
rect 29183 456 29239 458
rect 29183 404 29185 456
rect 29185 404 29237 456
rect 29237 404 29239 456
rect 29183 402 29239 404
rect 30431 456 30487 458
rect 30431 404 30433 456
rect 30433 404 30485 456
rect 30485 404 30487 456
rect 30431 402 30487 404
rect 31679 456 31735 458
rect 31679 404 31681 456
rect 31681 404 31733 456
rect 31733 404 31735 456
rect 31679 402 31735 404
rect 32927 456 32983 458
rect 32927 404 32929 456
rect 32929 404 32981 456
rect 32981 404 32983 456
rect 32927 402 32983 404
rect 34175 456 34231 458
rect 34175 404 34177 456
rect 34177 404 34229 456
rect 34229 404 34231 456
rect 34175 402 34231 404
rect 35423 456 35479 458
rect 35423 404 35425 456
rect 35425 404 35477 456
rect 35477 404 35479 456
rect 35423 402 35479 404
rect 36671 456 36727 458
rect 36671 404 36673 456
rect 36673 404 36725 456
rect 36725 404 36727 456
rect 36671 402 36727 404
rect 37919 456 37975 458
rect 37919 404 37921 456
rect 37921 404 37973 456
rect 37973 404 37975 456
rect 37919 402 37975 404
rect 39167 456 39223 458
rect 39167 404 39169 456
rect 39169 404 39221 456
rect 39221 404 39223 456
rect 39167 402 39223 404
rect 40415 456 40471 458
rect 40415 404 40417 456
rect 40417 404 40469 456
rect 40469 404 40471 456
rect 40415 402 40471 404
rect 1727 134 1783 136
rect 1727 82 1729 134
rect 1729 82 1781 134
rect 1781 82 1783 134
rect 1727 80 1783 82
rect 2975 134 3031 136
rect 2975 82 2977 134
rect 2977 82 3029 134
rect 3029 82 3031 134
rect 2975 80 3031 82
rect 4223 134 4279 136
rect 4223 82 4225 134
rect 4225 82 4277 134
rect 4277 82 4279 134
rect 4223 80 4279 82
rect 5471 134 5527 136
rect 5471 82 5473 134
rect 5473 82 5525 134
rect 5525 82 5527 134
rect 5471 80 5527 82
rect 6719 134 6775 136
rect 6719 82 6721 134
rect 6721 82 6773 134
rect 6773 82 6775 134
rect 6719 80 6775 82
rect 7967 134 8023 136
rect 7967 82 7969 134
rect 7969 82 8021 134
rect 8021 82 8023 134
rect 7967 80 8023 82
rect 9215 134 9271 136
rect 9215 82 9217 134
rect 9217 82 9269 134
rect 9269 82 9271 134
rect 9215 80 9271 82
rect 10463 134 10519 136
rect 10463 82 10465 134
rect 10465 82 10517 134
rect 10517 82 10519 134
rect 10463 80 10519 82
rect 11711 134 11767 136
rect 11711 82 11713 134
rect 11713 82 11765 134
rect 11765 82 11767 134
rect 11711 80 11767 82
rect 12959 134 13015 136
rect 12959 82 12961 134
rect 12961 82 13013 134
rect 13013 82 13015 134
rect 12959 80 13015 82
rect 14207 134 14263 136
rect 14207 82 14209 134
rect 14209 82 14261 134
rect 14261 82 14263 134
rect 14207 80 14263 82
rect 15455 134 15511 136
rect 15455 82 15457 134
rect 15457 82 15509 134
rect 15509 82 15511 134
rect 15455 80 15511 82
rect 16703 134 16759 136
rect 16703 82 16705 134
rect 16705 82 16757 134
rect 16757 82 16759 134
rect 16703 80 16759 82
rect 17951 134 18007 136
rect 17951 82 17953 134
rect 17953 82 18005 134
rect 18005 82 18007 134
rect 17951 80 18007 82
rect 19199 134 19255 136
rect 19199 82 19201 134
rect 19201 82 19253 134
rect 19253 82 19255 134
rect 19199 80 19255 82
rect 20447 134 20503 136
rect 20447 82 20449 134
rect 20449 82 20501 134
rect 20501 82 20503 134
rect 20447 80 20503 82
rect 21695 134 21751 136
rect 21695 82 21697 134
rect 21697 82 21749 134
rect 21749 82 21751 134
rect 21695 80 21751 82
rect 22943 134 22999 136
rect 22943 82 22945 134
rect 22945 82 22997 134
rect 22997 82 22999 134
rect 22943 80 22999 82
rect 24191 134 24247 136
rect 24191 82 24193 134
rect 24193 82 24245 134
rect 24245 82 24247 134
rect 24191 80 24247 82
rect 25439 134 25495 136
rect 25439 82 25441 134
rect 25441 82 25493 134
rect 25493 82 25495 134
rect 25439 80 25495 82
rect 26687 134 26743 136
rect 26687 82 26689 134
rect 26689 82 26741 134
rect 26741 82 26743 134
rect 26687 80 26743 82
rect 27935 134 27991 136
rect 27935 82 27937 134
rect 27937 82 27989 134
rect 27989 82 27991 134
rect 27935 80 27991 82
rect 29183 134 29239 136
rect 29183 82 29185 134
rect 29185 82 29237 134
rect 29237 82 29239 134
rect 29183 80 29239 82
rect 30431 134 30487 136
rect 30431 82 30433 134
rect 30433 82 30485 134
rect 30485 82 30487 134
rect 30431 80 30487 82
rect 31679 134 31735 136
rect 31679 82 31681 134
rect 31681 82 31733 134
rect 31733 82 31735 134
rect 31679 80 31735 82
rect 32927 134 32983 136
rect 32927 82 32929 134
rect 32929 82 32981 134
rect 32981 82 32983 134
rect 32927 80 32983 82
rect 34175 134 34231 136
rect 34175 82 34177 134
rect 34177 82 34229 134
rect 34229 82 34231 134
rect 34175 80 34231 82
rect 35423 134 35479 136
rect 35423 82 35425 134
rect 35425 82 35477 134
rect 35477 82 35479 134
rect 35423 80 35479 82
rect 36671 134 36727 136
rect 36671 82 36673 134
rect 36673 82 36725 134
rect 36725 82 36727 134
rect 36671 80 36727 82
rect 37919 134 37975 136
rect 37919 82 37921 134
rect 37921 82 37973 134
rect 37973 82 37975 134
rect 37919 80 37975 82
rect 39167 134 39223 136
rect 39167 82 39169 134
rect 39169 82 39221 134
rect 39221 82 39223 134
rect 39167 80 39223 82
rect 40415 134 40471 136
rect 40415 82 40417 134
rect 40417 82 40469 134
rect 40469 82 40471 134
rect 40415 80 40471 82
<< metal3 >>
rect 1464 2224 1530 2227
rect 2712 2224 2778 2227
rect 3960 2224 4026 2227
rect 5208 2224 5274 2227
rect 6456 2224 6522 2227
rect 7704 2224 7770 2227
rect 8952 2224 9018 2227
rect 10200 2224 10266 2227
rect 11448 2224 11514 2227
rect 12696 2224 12762 2227
rect 13944 2224 14010 2227
rect 15192 2224 15258 2227
rect 16440 2224 16506 2227
rect 17688 2224 17754 2227
rect 18936 2224 19002 2227
rect 20184 2224 20250 2227
rect 21432 2224 21498 2227
rect 22680 2224 22746 2227
rect 23928 2224 23994 2227
rect 25176 2224 25242 2227
rect 26424 2224 26490 2227
rect 27672 2224 27738 2227
rect 28920 2224 28986 2227
rect 30168 2224 30234 2227
rect 31416 2224 31482 2227
rect 32664 2224 32730 2227
rect 33912 2224 33978 2227
rect 35160 2224 35226 2227
rect 36408 2224 36474 2227
rect 37656 2224 37722 2227
rect 38904 2224 38970 2227
rect 40152 2224 40218 2227
rect 0 2222 40562 2224
rect 0 2166 1469 2222
rect 1525 2166 2717 2222
rect 2773 2166 3965 2222
rect 4021 2166 5213 2222
rect 5269 2166 6461 2222
rect 6517 2166 7709 2222
rect 7765 2166 8957 2222
rect 9013 2166 10205 2222
rect 10261 2166 11453 2222
rect 11509 2166 12701 2222
rect 12757 2166 13949 2222
rect 14005 2166 15197 2222
rect 15253 2166 16445 2222
rect 16501 2166 17693 2222
rect 17749 2166 18941 2222
rect 18997 2166 20189 2222
rect 20245 2166 21437 2222
rect 21493 2166 22685 2222
rect 22741 2166 23933 2222
rect 23989 2166 25181 2222
rect 25237 2166 26429 2222
rect 26485 2166 27677 2222
rect 27733 2166 28925 2222
rect 28981 2166 30173 2222
rect 30229 2166 31421 2222
rect 31477 2166 32669 2222
rect 32725 2166 33917 2222
rect 33973 2166 35165 2222
rect 35221 2166 36413 2222
rect 36469 2166 37661 2222
rect 37717 2166 38909 2222
rect 38965 2166 40157 2222
rect 40213 2166 40562 2222
rect 0 2164 40562 2166
rect 1464 2161 1530 2164
rect 2712 2161 2778 2164
rect 3960 2161 4026 2164
rect 5208 2161 5274 2164
rect 6456 2161 6522 2164
rect 7704 2161 7770 2164
rect 8952 2161 9018 2164
rect 10200 2161 10266 2164
rect 11448 2161 11514 2164
rect 12696 2161 12762 2164
rect 13944 2161 14010 2164
rect 15192 2161 15258 2164
rect 16440 2161 16506 2164
rect 17688 2161 17754 2164
rect 18936 2161 19002 2164
rect 20184 2161 20250 2164
rect 21432 2161 21498 2164
rect 22680 2161 22746 2164
rect 23928 2161 23994 2164
rect 25176 2161 25242 2164
rect 26424 2161 26490 2164
rect 27672 2161 27738 2164
rect 28920 2161 28986 2164
rect 30168 2161 30234 2164
rect 31416 2161 31482 2164
rect 32664 2161 32730 2164
rect 33912 2161 33978 2164
rect 35160 2161 35226 2164
rect 36408 2161 36474 2164
rect 37656 2161 37722 2164
rect 38904 2161 38970 2164
rect 40152 2161 40218 2164
rect 1776 2070 1874 2091
rect 1776 2014 1797 2070
rect 1853 2014 1874 2070
rect 1776 1993 1874 2014
rect 3024 2070 3122 2091
rect 3024 2014 3045 2070
rect 3101 2014 3122 2070
rect 3024 1993 3122 2014
rect 4272 2070 4370 2091
rect 4272 2014 4293 2070
rect 4349 2014 4370 2070
rect 4272 1993 4370 2014
rect 5520 2070 5618 2091
rect 5520 2014 5541 2070
rect 5597 2014 5618 2070
rect 5520 1993 5618 2014
rect 6768 2070 6866 2091
rect 6768 2014 6789 2070
rect 6845 2014 6866 2070
rect 6768 1993 6866 2014
rect 8016 2070 8114 2091
rect 8016 2014 8037 2070
rect 8093 2014 8114 2070
rect 8016 1993 8114 2014
rect 9264 2070 9362 2091
rect 9264 2014 9285 2070
rect 9341 2014 9362 2070
rect 9264 1993 9362 2014
rect 10512 2070 10610 2091
rect 10512 2014 10533 2070
rect 10589 2014 10610 2070
rect 10512 1993 10610 2014
rect 11760 2070 11858 2091
rect 11760 2014 11781 2070
rect 11837 2014 11858 2070
rect 11760 1993 11858 2014
rect 13008 2070 13106 2091
rect 13008 2014 13029 2070
rect 13085 2014 13106 2070
rect 13008 1993 13106 2014
rect 14256 2070 14354 2091
rect 14256 2014 14277 2070
rect 14333 2014 14354 2070
rect 14256 1993 14354 2014
rect 15504 2070 15602 2091
rect 15504 2014 15525 2070
rect 15581 2014 15602 2070
rect 15504 1993 15602 2014
rect 16752 2070 16850 2091
rect 16752 2014 16773 2070
rect 16829 2014 16850 2070
rect 16752 1993 16850 2014
rect 18000 2070 18098 2091
rect 18000 2014 18021 2070
rect 18077 2014 18098 2070
rect 18000 1993 18098 2014
rect 19248 2070 19346 2091
rect 19248 2014 19269 2070
rect 19325 2014 19346 2070
rect 19248 1993 19346 2014
rect 20496 2070 20594 2091
rect 20496 2014 20517 2070
rect 20573 2014 20594 2070
rect 20496 1993 20594 2014
rect 21744 2070 21842 2091
rect 21744 2014 21765 2070
rect 21821 2014 21842 2070
rect 21744 1993 21842 2014
rect 22992 2070 23090 2091
rect 22992 2014 23013 2070
rect 23069 2014 23090 2070
rect 22992 1993 23090 2014
rect 24240 2070 24338 2091
rect 24240 2014 24261 2070
rect 24317 2014 24338 2070
rect 24240 1993 24338 2014
rect 25488 2070 25586 2091
rect 25488 2014 25509 2070
rect 25565 2014 25586 2070
rect 25488 1993 25586 2014
rect 26736 2070 26834 2091
rect 26736 2014 26757 2070
rect 26813 2014 26834 2070
rect 26736 1993 26834 2014
rect 27984 2070 28082 2091
rect 27984 2014 28005 2070
rect 28061 2014 28082 2070
rect 27984 1993 28082 2014
rect 29232 2070 29330 2091
rect 29232 2014 29253 2070
rect 29309 2014 29330 2070
rect 29232 1993 29330 2014
rect 30480 2070 30578 2091
rect 30480 2014 30501 2070
rect 30557 2014 30578 2070
rect 30480 1993 30578 2014
rect 31728 2070 31826 2091
rect 31728 2014 31749 2070
rect 31805 2014 31826 2070
rect 31728 1993 31826 2014
rect 32976 2070 33074 2091
rect 32976 2014 32997 2070
rect 33053 2014 33074 2070
rect 32976 1993 33074 2014
rect 34224 2070 34322 2091
rect 34224 2014 34245 2070
rect 34301 2014 34322 2070
rect 34224 1993 34322 2014
rect 35472 2070 35570 2091
rect 35472 2014 35493 2070
rect 35549 2014 35570 2070
rect 35472 1993 35570 2014
rect 36720 2070 36818 2091
rect 36720 2014 36741 2070
rect 36797 2014 36818 2070
rect 36720 1993 36818 2014
rect 37968 2070 38066 2091
rect 37968 2014 37989 2070
rect 38045 2014 38066 2070
rect 37968 1993 38066 2014
rect 39216 2070 39314 2091
rect 39216 2014 39237 2070
rect 39293 2014 39314 2070
rect 39216 1993 39314 2014
rect 40464 2070 40562 2091
rect 40464 2014 40485 2070
rect 40541 2014 40562 2070
rect 40464 1993 40562 2014
rect 1694 1296 1792 1317
rect 1694 1240 1715 1296
rect 1771 1240 1792 1296
rect 1694 1219 1792 1240
rect 2942 1296 3040 1317
rect 2942 1240 2963 1296
rect 3019 1240 3040 1296
rect 2942 1219 3040 1240
rect 4190 1296 4288 1317
rect 4190 1240 4211 1296
rect 4267 1240 4288 1296
rect 4190 1219 4288 1240
rect 5438 1296 5536 1317
rect 5438 1240 5459 1296
rect 5515 1240 5536 1296
rect 5438 1219 5536 1240
rect 6686 1296 6784 1317
rect 6686 1240 6707 1296
rect 6763 1240 6784 1296
rect 6686 1219 6784 1240
rect 7934 1296 8032 1317
rect 7934 1240 7955 1296
rect 8011 1240 8032 1296
rect 7934 1219 8032 1240
rect 9182 1296 9280 1317
rect 9182 1240 9203 1296
rect 9259 1240 9280 1296
rect 9182 1219 9280 1240
rect 10430 1296 10528 1317
rect 10430 1240 10451 1296
rect 10507 1240 10528 1296
rect 10430 1219 10528 1240
rect 11678 1296 11776 1317
rect 11678 1240 11699 1296
rect 11755 1240 11776 1296
rect 11678 1219 11776 1240
rect 12926 1296 13024 1317
rect 12926 1240 12947 1296
rect 13003 1240 13024 1296
rect 12926 1219 13024 1240
rect 14174 1296 14272 1317
rect 14174 1240 14195 1296
rect 14251 1240 14272 1296
rect 14174 1219 14272 1240
rect 15422 1296 15520 1317
rect 15422 1240 15443 1296
rect 15499 1240 15520 1296
rect 15422 1219 15520 1240
rect 16670 1296 16768 1317
rect 16670 1240 16691 1296
rect 16747 1240 16768 1296
rect 16670 1219 16768 1240
rect 17918 1296 18016 1317
rect 17918 1240 17939 1296
rect 17995 1240 18016 1296
rect 17918 1219 18016 1240
rect 19166 1296 19264 1317
rect 19166 1240 19187 1296
rect 19243 1240 19264 1296
rect 19166 1219 19264 1240
rect 20414 1296 20512 1317
rect 20414 1240 20435 1296
rect 20491 1240 20512 1296
rect 20414 1219 20512 1240
rect 21662 1296 21760 1317
rect 21662 1240 21683 1296
rect 21739 1240 21760 1296
rect 21662 1219 21760 1240
rect 22910 1296 23008 1317
rect 22910 1240 22931 1296
rect 22987 1240 23008 1296
rect 22910 1219 23008 1240
rect 24158 1296 24256 1317
rect 24158 1240 24179 1296
rect 24235 1240 24256 1296
rect 24158 1219 24256 1240
rect 25406 1296 25504 1317
rect 25406 1240 25427 1296
rect 25483 1240 25504 1296
rect 25406 1219 25504 1240
rect 26654 1296 26752 1317
rect 26654 1240 26675 1296
rect 26731 1240 26752 1296
rect 26654 1219 26752 1240
rect 27902 1296 28000 1317
rect 27902 1240 27923 1296
rect 27979 1240 28000 1296
rect 27902 1219 28000 1240
rect 29150 1296 29248 1317
rect 29150 1240 29171 1296
rect 29227 1240 29248 1296
rect 29150 1219 29248 1240
rect 30398 1296 30496 1317
rect 30398 1240 30419 1296
rect 30475 1240 30496 1296
rect 30398 1219 30496 1240
rect 31646 1296 31744 1317
rect 31646 1240 31667 1296
rect 31723 1240 31744 1296
rect 31646 1219 31744 1240
rect 32894 1296 32992 1317
rect 32894 1240 32915 1296
rect 32971 1240 32992 1296
rect 32894 1219 32992 1240
rect 34142 1296 34240 1317
rect 34142 1240 34163 1296
rect 34219 1240 34240 1296
rect 34142 1219 34240 1240
rect 35390 1296 35488 1317
rect 35390 1240 35411 1296
rect 35467 1240 35488 1296
rect 35390 1219 35488 1240
rect 36638 1296 36736 1317
rect 36638 1240 36659 1296
rect 36715 1240 36736 1296
rect 36638 1219 36736 1240
rect 37886 1296 37984 1317
rect 37886 1240 37907 1296
rect 37963 1240 37984 1296
rect 37886 1219 37984 1240
rect 39134 1296 39232 1317
rect 39134 1240 39155 1296
rect 39211 1240 39232 1296
rect 39134 1219 39232 1240
rect 40382 1296 40480 1317
rect 40382 1240 40403 1296
rect 40459 1240 40480 1296
rect 40382 1219 40480 1240
rect 1706 458 1804 479
rect 1706 402 1727 458
rect 1783 402 1804 458
rect 1706 381 1804 402
rect 2954 458 3052 479
rect 2954 402 2975 458
rect 3031 402 3052 458
rect 2954 381 3052 402
rect 4202 458 4300 479
rect 4202 402 4223 458
rect 4279 402 4300 458
rect 4202 381 4300 402
rect 5450 458 5548 479
rect 5450 402 5471 458
rect 5527 402 5548 458
rect 5450 381 5548 402
rect 6698 458 6796 479
rect 6698 402 6719 458
rect 6775 402 6796 458
rect 6698 381 6796 402
rect 7946 458 8044 479
rect 7946 402 7967 458
rect 8023 402 8044 458
rect 7946 381 8044 402
rect 9194 458 9292 479
rect 9194 402 9215 458
rect 9271 402 9292 458
rect 9194 381 9292 402
rect 10442 458 10540 479
rect 10442 402 10463 458
rect 10519 402 10540 458
rect 10442 381 10540 402
rect 11690 458 11788 479
rect 11690 402 11711 458
rect 11767 402 11788 458
rect 11690 381 11788 402
rect 12938 458 13036 479
rect 12938 402 12959 458
rect 13015 402 13036 458
rect 12938 381 13036 402
rect 14186 458 14284 479
rect 14186 402 14207 458
rect 14263 402 14284 458
rect 14186 381 14284 402
rect 15434 458 15532 479
rect 15434 402 15455 458
rect 15511 402 15532 458
rect 15434 381 15532 402
rect 16682 458 16780 479
rect 16682 402 16703 458
rect 16759 402 16780 458
rect 16682 381 16780 402
rect 17930 458 18028 479
rect 17930 402 17951 458
rect 18007 402 18028 458
rect 17930 381 18028 402
rect 19178 458 19276 479
rect 19178 402 19199 458
rect 19255 402 19276 458
rect 19178 381 19276 402
rect 20426 458 20524 479
rect 20426 402 20447 458
rect 20503 402 20524 458
rect 20426 381 20524 402
rect 21674 458 21772 479
rect 21674 402 21695 458
rect 21751 402 21772 458
rect 21674 381 21772 402
rect 22922 458 23020 479
rect 22922 402 22943 458
rect 22999 402 23020 458
rect 22922 381 23020 402
rect 24170 458 24268 479
rect 24170 402 24191 458
rect 24247 402 24268 458
rect 24170 381 24268 402
rect 25418 458 25516 479
rect 25418 402 25439 458
rect 25495 402 25516 458
rect 25418 381 25516 402
rect 26666 458 26764 479
rect 26666 402 26687 458
rect 26743 402 26764 458
rect 26666 381 26764 402
rect 27914 458 28012 479
rect 27914 402 27935 458
rect 27991 402 28012 458
rect 27914 381 28012 402
rect 29162 458 29260 479
rect 29162 402 29183 458
rect 29239 402 29260 458
rect 29162 381 29260 402
rect 30410 458 30508 479
rect 30410 402 30431 458
rect 30487 402 30508 458
rect 30410 381 30508 402
rect 31658 458 31756 479
rect 31658 402 31679 458
rect 31735 402 31756 458
rect 31658 381 31756 402
rect 32906 458 33004 479
rect 32906 402 32927 458
rect 32983 402 33004 458
rect 32906 381 33004 402
rect 34154 458 34252 479
rect 34154 402 34175 458
rect 34231 402 34252 458
rect 34154 381 34252 402
rect 35402 458 35500 479
rect 35402 402 35423 458
rect 35479 402 35500 458
rect 35402 381 35500 402
rect 36650 458 36748 479
rect 36650 402 36671 458
rect 36727 402 36748 458
rect 36650 381 36748 402
rect 37898 458 37996 479
rect 37898 402 37919 458
rect 37975 402 37996 458
rect 37898 381 37996 402
rect 39146 458 39244 479
rect 39146 402 39167 458
rect 39223 402 39244 458
rect 39146 381 39244 402
rect 40394 458 40492 479
rect 40394 402 40415 458
rect 40471 402 40492 458
rect 40394 381 40492 402
rect 1706 136 1804 157
rect 1706 80 1727 136
rect 1783 80 1804 136
rect 1706 59 1804 80
rect 2954 136 3052 157
rect 2954 80 2975 136
rect 3031 80 3052 136
rect 2954 59 3052 80
rect 4202 136 4300 157
rect 4202 80 4223 136
rect 4279 80 4300 136
rect 4202 59 4300 80
rect 5450 136 5548 157
rect 5450 80 5471 136
rect 5527 80 5548 136
rect 5450 59 5548 80
rect 6698 136 6796 157
rect 6698 80 6719 136
rect 6775 80 6796 136
rect 6698 59 6796 80
rect 7946 136 8044 157
rect 7946 80 7967 136
rect 8023 80 8044 136
rect 7946 59 8044 80
rect 9194 136 9292 157
rect 9194 80 9215 136
rect 9271 80 9292 136
rect 9194 59 9292 80
rect 10442 136 10540 157
rect 10442 80 10463 136
rect 10519 80 10540 136
rect 10442 59 10540 80
rect 11690 136 11788 157
rect 11690 80 11711 136
rect 11767 80 11788 136
rect 11690 59 11788 80
rect 12938 136 13036 157
rect 12938 80 12959 136
rect 13015 80 13036 136
rect 12938 59 13036 80
rect 14186 136 14284 157
rect 14186 80 14207 136
rect 14263 80 14284 136
rect 14186 59 14284 80
rect 15434 136 15532 157
rect 15434 80 15455 136
rect 15511 80 15532 136
rect 15434 59 15532 80
rect 16682 136 16780 157
rect 16682 80 16703 136
rect 16759 80 16780 136
rect 16682 59 16780 80
rect 17930 136 18028 157
rect 17930 80 17951 136
rect 18007 80 18028 136
rect 17930 59 18028 80
rect 19178 136 19276 157
rect 19178 80 19199 136
rect 19255 80 19276 136
rect 19178 59 19276 80
rect 20426 136 20524 157
rect 20426 80 20447 136
rect 20503 80 20524 136
rect 20426 59 20524 80
rect 21674 136 21772 157
rect 21674 80 21695 136
rect 21751 80 21772 136
rect 21674 59 21772 80
rect 22922 136 23020 157
rect 22922 80 22943 136
rect 22999 80 23020 136
rect 22922 59 23020 80
rect 24170 136 24268 157
rect 24170 80 24191 136
rect 24247 80 24268 136
rect 24170 59 24268 80
rect 25418 136 25516 157
rect 25418 80 25439 136
rect 25495 80 25516 136
rect 25418 59 25516 80
rect 26666 136 26764 157
rect 26666 80 26687 136
rect 26743 80 26764 136
rect 26666 59 26764 80
rect 27914 136 28012 157
rect 27914 80 27935 136
rect 27991 80 28012 136
rect 27914 59 28012 80
rect 29162 136 29260 157
rect 29162 80 29183 136
rect 29239 80 29260 136
rect 29162 59 29260 80
rect 30410 136 30508 157
rect 30410 80 30431 136
rect 30487 80 30508 136
rect 30410 59 30508 80
rect 31658 136 31756 157
rect 31658 80 31679 136
rect 31735 80 31756 136
rect 31658 59 31756 80
rect 32906 136 33004 157
rect 32906 80 32927 136
rect 32983 80 33004 136
rect 32906 59 33004 80
rect 34154 136 34252 157
rect 34154 80 34175 136
rect 34231 80 34252 136
rect 34154 59 34252 80
rect 35402 136 35500 157
rect 35402 80 35423 136
rect 35479 80 35500 136
rect 35402 59 35500 80
rect 36650 136 36748 157
rect 36650 80 36671 136
rect 36727 80 36748 136
rect 36650 59 36748 80
rect 37898 136 37996 157
rect 37898 80 37919 136
rect 37975 80 37996 136
rect 37898 59 37996 80
rect 39146 136 39244 157
rect 39146 80 39167 136
rect 39223 80 39244 136
rect 39146 59 39244 80
rect 40394 136 40492 157
rect 40394 80 40415 136
rect 40471 80 40492 136
rect 40394 59 40492 80
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_0
timestamp 1666464484
transform 1 0 2622 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_1
timestamp 1666464484
transform 1 0 1374 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_2
timestamp 1666464484
transform 1 0 8862 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_3
timestamp 1666464484
transform 1 0 7614 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_4
timestamp 1666464484
transform 1 0 6366 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_5
timestamp 1666464484
transform 1 0 5118 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_6
timestamp 1666464484
transform 1 0 3870 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_7
timestamp 1666464484
transform 1 0 18846 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_8
timestamp 1666464484
transform 1 0 17598 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_9
timestamp 1666464484
transform 1 0 16350 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_10
timestamp 1666464484
transform 1 0 15102 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_11
timestamp 1666464484
transform 1 0 13854 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_12
timestamp 1666464484
transform 1 0 12606 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_13
timestamp 1666464484
transform 1 0 11358 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_14
timestamp 1666464484
transform 1 0 10110 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_15
timestamp 1666464484
transform 1 0 25086 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_16
timestamp 1666464484
transform 1 0 23838 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_17
timestamp 1666464484
transform 1 0 22590 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_18
timestamp 1666464484
transform 1 0 28830 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_19
timestamp 1666464484
transform 1 0 27582 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_20
timestamp 1666464484
transform 1 0 26334 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_21
timestamp 1666464484
transform 1 0 40062 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_22
timestamp 1666464484
transform 1 0 38814 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_23
timestamp 1666464484
transform 1 0 37566 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_24
timestamp 1666464484
transform 1 0 36318 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_25
timestamp 1666464484
transform 1 0 35070 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_26
timestamp 1666464484
transform 1 0 33822 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_27
timestamp 1666464484
transform 1 0 32574 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_28
timestamp 1666464484
transform 1 0 31326 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_29
timestamp 1666464484
transform 1 0 30078 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_30
timestamp 1666464484
transform 1 0 21342 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_31
timestamp 1666464484
transform 1 0 20094 0 1 0
box -541 0 937 2256
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_0
timestamp 1666464484
transform 1 0 1792 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_1
timestamp 1666464484
transform 1 0 5466 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_2
timestamp 1666464484
transform 1 0 5536 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_3
timestamp 1666464484
transform 1 0 4218 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_4
timestamp 1666464484
transform 1 0 4206 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_5
timestamp 1666464484
transform 1 0 4218 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_6
timestamp 1666464484
transform 1 0 4288 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_7
timestamp 1666464484
transform 1 0 2970 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_8
timestamp 1666464484
transform 1 0 2958 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_9
timestamp 1666464484
transform 1 0 2970 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_10
timestamp 1666464484
transform 1 0 3040 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_11
timestamp 1666464484
transform 1 0 1722 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_12
timestamp 1666464484
transform 1 0 1710 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_13
timestamp 1666464484
transform 1 0 1722 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_14
timestamp 1666464484
transform 1 0 10458 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_15
timestamp 1666464484
transform 1 0 10446 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_16
timestamp 1666464484
transform 1 0 10458 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_17
timestamp 1666464484
transform 1 0 10528 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_18
timestamp 1666464484
transform 1 0 9210 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_19
timestamp 1666464484
transform 1 0 9198 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_20
timestamp 1666464484
transform 1 0 9210 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_21
timestamp 1666464484
transform 1 0 10200 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_22
timestamp 1666464484
transform 1 0 8952 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_23
timestamp 1666464484
transform 1 0 7704 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_24
timestamp 1666464484
transform 1 0 6456 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_25
timestamp 1666464484
transform 1 0 5208 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_26
timestamp 1666464484
transform 1 0 3960 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_27
timestamp 1666464484
transform 1 0 2712 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_28
timestamp 1666464484
transform 1 0 1464 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_29
timestamp 1666464484
transform 1 0 9280 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_30
timestamp 1666464484
transform 1 0 7962 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_31
timestamp 1666464484
transform 1 0 7950 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_32
timestamp 1666464484
transform 1 0 7962 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_33
timestamp 1666464484
transform 1 0 8032 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_34
timestamp 1666464484
transform 1 0 6714 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_35
timestamp 1666464484
transform 1 0 6702 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_36
timestamp 1666464484
transform 1 0 6714 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_37
timestamp 1666464484
transform 1 0 6784 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_38
timestamp 1666464484
transform 1 0 5466 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_39
timestamp 1666464484
transform 1 0 5454 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_40
timestamp 1666464484
transform 1 0 11776 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_41
timestamp 1666464484
transform 1 0 20442 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_42
timestamp 1666464484
transform 1 0 20430 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_43
timestamp 1666464484
transform 1 0 20442 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_44
timestamp 1666464484
transform 1 0 20512 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_45
timestamp 1666464484
transform 1 0 19194 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_46
timestamp 1666464484
transform 1 0 19182 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_47
timestamp 1666464484
transform 1 0 19194 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_48
timestamp 1666464484
transform 1 0 19264 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_49
timestamp 1666464484
transform 1 0 20184 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_50
timestamp 1666464484
transform 1 0 18936 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_51
timestamp 1666464484
transform 1 0 17688 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_52
timestamp 1666464484
transform 1 0 16440 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_53
timestamp 1666464484
transform 1 0 15192 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_54
timestamp 1666464484
transform 1 0 13944 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_55
timestamp 1666464484
transform 1 0 12696 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_56
timestamp 1666464484
transform 1 0 11448 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_57
timestamp 1666464484
transform 1 0 17946 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_58
timestamp 1666464484
transform 1 0 17934 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_59
timestamp 1666464484
transform 1 0 17946 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_60
timestamp 1666464484
transform 1 0 18016 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_61
timestamp 1666464484
transform 1 0 16698 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_62
timestamp 1666464484
transform 1 0 16686 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_63
timestamp 1666464484
transform 1 0 16698 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_64
timestamp 1666464484
transform 1 0 16768 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_65
timestamp 1666464484
transform 1 0 15450 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_66
timestamp 1666464484
transform 1 0 15438 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_67
timestamp 1666464484
transform 1 0 15450 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_68
timestamp 1666464484
transform 1 0 15520 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_69
timestamp 1666464484
transform 1 0 14202 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_70
timestamp 1666464484
transform 1 0 14190 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_71
timestamp 1666464484
transform 1 0 14202 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_72
timestamp 1666464484
transform 1 0 14272 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_73
timestamp 1666464484
transform 1 0 12954 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_74
timestamp 1666464484
transform 1 0 12942 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_75
timestamp 1666464484
transform 1 0 12954 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_76
timestamp 1666464484
transform 1 0 13024 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_77
timestamp 1666464484
transform 1 0 11706 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_78
timestamp 1666464484
transform 1 0 11694 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_79
timestamp 1666464484
transform 1 0 11706 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_80
timestamp 1666464484
transform 1 0 21690 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_81
timestamp 1666464484
transform 1 0 21760 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_82
timestamp 1666464484
transform 1 0 30426 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_83
timestamp 1666464484
transform 1 0 30414 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_84
timestamp 1666464484
transform 1 0 30426 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_85
timestamp 1666464484
transform 1 0 30168 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_86
timestamp 1666464484
transform 1 0 28920 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_87
timestamp 1666464484
transform 1 0 27672 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_88
timestamp 1666464484
transform 1 0 26424 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_89
timestamp 1666464484
transform 1 0 25176 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_90
timestamp 1666464484
transform 1 0 23928 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_91
timestamp 1666464484
transform 1 0 22680 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_92
timestamp 1666464484
transform 1 0 21432 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_93
timestamp 1666464484
transform 1 0 30496 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_94
timestamp 1666464484
transform 1 0 29178 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_95
timestamp 1666464484
transform 1 0 29166 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_96
timestamp 1666464484
transform 1 0 29178 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_97
timestamp 1666464484
transform 1 0 29248 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_98
timestamp 1666464484
transform 1 0 27930 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_99
timestamp 1666464484
transform 1 0 27918 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_100
timestamp 1666464484
transform 1 0 27930 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_101
timestamp 1666464484
transform 1 0 28000 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_102
timestamp 1666464484
transform 1 0 26682 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_103
timestamp 1666464484
transform 1 0 26670 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_104
timestamp 1666464484
transform 1 0 26682 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_105
timestamp 1666464484
transform 1 0 26752 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_106
timestamp 1666464484
transform 1 0 25434 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_107
timestamp 1666464484
transform 1 0 25422 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_108
timestamp 1666464484
transform 1 0 25434 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_109
timestamp 1666464484
transform 1 0 25504 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_110
timestamp 1666464484
transform 1 0 24186 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_111
timestamp 1666464484
transform 1 0 24174 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_112
timestamp 1666464484
transform 1 0 24186 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_113
timestamp 1666464484
transform 1 0 24256 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_114
timestamp 1666464484
transform 1 0 22938 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_115
timestamp 1666464484
transform 1 0 22926 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_116
timestamp 1666464484
transform 1 0 22938 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_117
timestamp 1666464484
transform 1 0 23008 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_118
timestamp 1666464484
transform 1 0 21690 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_119
timestamp 1666464484
transform 1 0 21678 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_120
timestamp 1666464484
transform 1 0 40152 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_121
timestamp 1666464484
transform 1 0 38904 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_122
timestamp 1666464484
transform 1 0 37656 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_123
timestamp 1666464484
transform 1 0 36408 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_124
timestamp 1666464484
transform 1 0 35160 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_125
timestamp 1666464484
transform 1 0 33912 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_126
timestamp 1666464484
transform 1 0 32664 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_127
timestamp 1666464484
transform 1 0 31416 0 1 2157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_128
timestamp 1666464484
transform 1 0 40410 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_129
timestamp 1666464484
transform 1 0 40398 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_130
timestamp 1666464484
transform 1 0 40410 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_131
timestamp 1666464484
transform 1 0 40480 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_132
timestamp 1666464484
transform 1 0 39162 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_133
timestamp 1666464484
transform 1 0 39150 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_134
timestamp 1666464484
transform 1 0 39162 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_135
timestamp 1666464484
transform 1 0 39232 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_136
timestamp 1666464484
transform 1 0 37914 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_137
timestamp 1666464484
transform 1 0 37902 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_138
timestamp 1666464484
transform 1 0 37914 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_139
timestamp 1666464484
transform 1 0 37984 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_140
timestamp 1666464484
transform 1 0 36666 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_141
timestamp 1666464484
transform 1 0 36654 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_142
timestamp 1666464484
transform 1 0 36666 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_143
timestamp 1666464484
transform 1 0 36736 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_144
timestamp 1666464484
transform 1 0 35418 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_145
timestamp 1666464484
transform 1 0 35406 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_146
timestamp 1666464484
transform 1 0 35418 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_147
timestamp 1666464484
transform 1 0 35488 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_148
timestamp 1666464484
transform 1 0 34170 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_149
timestamp 1666464484
transform 1 0 34158 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_150
timestamp 1666464484
transform 1 0 34170 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_151
timestamp 1666464484
transform 1 0 34240 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_152
timestamp 1666464484
transform 1 0 32922 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_153
timestamp 1666464484
transform 1 0 32910 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_154
timestamp 1666464484
transform 1 0 32922 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_155
timestamp 1666464484
transform 1 0 32992 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_156
timestamp 1666464484
transform 1 0 31674 0 1 393
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_157
timestamp 1666464484
transform 1 0 31662 0 1 1231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_158
timestamp 1666464484
transform 1 0 31674 0 1 71
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_159
timestamp 1666464484
transform 1 0 31744 0 1 2005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1666464484
transform 1 0 1793 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1666464484
transform 1 0 5467 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1666464484
transform 1 0 5537 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_3
timestamp 1666464484
transform 1 0 4219 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_4
timestamp 1666464484
transform 1 0 4207 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_5
timestamp 1666464484
transform 1 0 4219 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_6
timestamp 1666464484
transform 1 0 4289 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_7
timestamp 1666464484
transform 1 0 2971 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_8
timestamp 1666464484
transform 1 0 2959 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_9
timestamp 1666464484
transform 1 0 2971 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_10
timestamp 1666464484
transform 1 0 3041 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_11
timestamp 1666464484
transform 1 0 1723 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_12
timestamp 1666464484
transform 1 0 1711 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_13
timestamp 1666464484
transform 1 0 1723 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_14
timestamp 1666464484
transform 1 0 10459 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_15
timestamp 1666464484
transform 1 0 10447 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_16
timestamp 1666464484
transform 1 0 10459 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_17
timestamp 1666464484
transform 1 0 10529 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_18
timestamp 1666464484
transform 1 0 9211 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_19
timestamp 1666464484
transform 1 0 9199 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_20
timestamp 1666464484
transform 1 0 10201 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_21
timestamp 1666464484
transform 1 0 8953 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_22
timestamp 1666464484
transform 1 0 7705 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_23
timestamp 1666464484
transform 1 0 6457 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_24
timestamp 1666464484
transform 1 0 5209 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_25
timestamp 1666464484
transform 1 0 3961 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_26
timestamp 1666464484
transform 1 0 2713 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_27
timestamp 1666464484
transform 1 0 1465 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_28
timestamp 1666464484
transform 1 0 9211 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_29
timestamp 1666464484
transform 1 0 9281 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_30
timestamp 1666464484
transform 1 0 7963 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_31
timestamp 1666464484
transform 1 0 7951 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_32
timestamp 1666464484
transform 1 0 7963 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_33
timestamp 1666464484
transform 1 0 8033 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_34
timestamp 1666464484
transform 1 0 6715 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_35
timestamp 1666464484
transform 1 0 6703 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_36
timestamp 1666464484
transform 1 0 6715 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_37
timestamp 1666464484
transform 1 0 6785 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_38
timestamp 1666464484
transform 1 0 5467 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_39
timestamp 1666464484
transform 1 0 5455 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_40
timestamp 1666464484
transform 1 0 11777 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_41
timestamp 1666464484
transform 1 0 20443 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_42
timestamp 1666464484
transform 1 0 20431 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_43
timestamp 1666464484
transform 1 0 20443 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_44
timestamp 1666464484
transform 1 0 20513 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_45
timestamp 1666464484
transform 1 0 19195 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_46
timestamp 1666464484
transform 1 0 19183 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_47
timestamp 1666464484
transform 1 0 19195 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_48
timestamp 1666464484
transform 1 0 20185 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_49
timestamp 1666464484
transform 1 0 18937 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_50
timestamp 1666464484
transform 1 0 17689 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_51
timestamp 1666464484
transform 1 0 16441 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_52
timestamp 1666464484
transform 1 0 15193 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_53
timestamp 1666464484
transform 1 0 13945 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_54
timestamp 1666464484
transform 1 0 12697 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_55
timestamp 1666464484
transform 1 0 11449 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_56
timestamp 1666464484
transform 1 0 19265 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_57
timestamp 1666464484
transform 1 0 17947 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_58
timestamp 1666464484
transform 1 0 17935 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_59
timestamp 1666464484
transform 1 0 17947 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_60
timestamp 1666464484
transform 1 0 18017 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_61
timestamp 1666464484
transform 1 0 16699 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_62
timestamp 1666464484
transform 1 0 16687 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_63
timestamp 1666464484
transform 1 0 16699 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_64
timestamp 1666464484
transform 1 0 16769 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_65
timestamp 1666464484
transform 1 0 15451 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_66
timestamp 1666464484
transform 1 0 15439 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_67
timestamp 1666464484
transform 1 0 15451 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_68
timestamp 1666464484
transform 1 0 15521 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_69
timestamp 1666464484
transform 1 0 14203 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_70
timestamp 1666464484
transform 1 0 14191 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_71
timestamp 1666464484
transform 1 0 14203 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_72
timestamp 1666464484
transform 1 0 14273 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_73
timestamp 1666464484
transform 1 0 12955 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_74
timestamp 1666464484
transform 1 0 12943 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_75
timestamp 1666464484
transform 1 0 12955 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_76
timestamp 1666464484
transform 1 0 13025 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_77
timestamp 1666464484
transform 1 0 11707 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_78
timestamp 1666464484
transform 1 0 11695 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_79
timestamp 1666464484
transform 1 0 11707 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_80
timestamp 1666464484
transform 1 0 21691 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_81
timestamp 1666464484
transform 1 0 21761 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_82
timestamp 1666464484
transform 1 0 30427 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_83
timestamp 1666464484
transform 1 0 30415 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_84
timestamp 1666464484
transform 1 0 30427 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_85
timestamp 1666464484
transform 1 0 30169 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_86
timestamp 1666464484
transform 1 0 28921 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_87
timestamp 1666464484
transform 1 0 27673 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_88
timestamp 1666464484
transform 1 0 26425 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_89
timestamp 1666464484
transform 1 0 25177 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_90
timestamp 1666464484
transform 1 0 23929 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_91
timestamp 1666464484
transform 1 0 22681 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_92
timestamp 1666464484
transform 1 0 21433 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_93
timestamp 1666464484
transform 1 0 30497 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_94
timestamp 1666464484
transform 1 0 29179 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_95
timestamp 1666464484
transform 1 0 29167 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_96
timestamp 1666464484
transform 1 0 29179 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_97
timestamp 1666464484
transform 1 0 29249 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_98
timestamp 1666464484
transform 1 0 27931 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_99
timestamp 1666464484
transform 1 0 27919 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_100
timestamp 1666464484
transform 1 0 27931 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_101
timestamp 1666464484
transform 1 0 28001 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_102
timestamp 1666464484
transform 1 0 26683 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_103
timestamp 1666464484
transform 1 0 26671 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_104
timestamp 1666464484
transform 1 0 26683 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_105
timestamp 1666464484
transform 1 0 26753 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_106
timestamp 1666464484
transform 1 0 25435 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_107
timestamp 1666464484
transform 1 0 25423 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_108
timestamp 1666464484
transform 1 0 25435 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_109
timestamp 1666464484
transform 1 0 25505 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_110
timestamp 1666464484
transform 1 0 24187 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_111
timestamp 1666464484
transform 1 0 24175 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_112
timestamp 1666464484
transform 1 0 24187 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_113
timestamp 1666464484
transform 1 0 24257 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_114
timestamp 1666464484
transform 1 0 22939 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_115
timestamp 1666464484
transform 1 0 22927 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_116
timestamp 1666464484
transform 1 0 22939 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_117
timestamp 1666464484
transform 1 0 23009 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_118
timestamp 1666464484
transform 1 0 21691 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_119
timestamp 1666464484
transform 1 0 21679 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_120
timestamp 1666464484
transform 1 0 40153 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_121
timestamp 1666464484
transform 1 0 38905 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_122
timestamp 1666464484
transform 1 0 37657 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_123
timestamp 1666464484
transform 1 0 36409 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_124
timestamp 1666464484
transform 1 0 35161 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_125
timestamp 1666464484
transform 1 0 33913 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_126
timestamp 1666464484
transform 1 0 32665 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_127
timestamp 1666464484
transform 1 0 31417 0 1 2162
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_128
timestamp 1666464484
transform 1 0 40411 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_129
timestamp 1666464484
transform 1 0 40399 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_130
timestamp 1666464484
transform 1 0 40411 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_131
timestamp 1666464484
transform 1 0 40481 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_132
timestamp 1666464484
transform 1 0 39163 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_133
timestamp 1666464484
transform 1 0 39151 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_134
timestamp 1666464484
transform 1 0 39163 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_135
timestamp 1666464484
transform 1 0 39233 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_136
timestamp 1666464484
transform 1 0 37915 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_137
timestamp 1666464484
transform 1 0 37903 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_138
timestamp 1666464484
transform 1 0 37915 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_139
timestamp 1666464484
transform 1 0 37985 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_140
timestamp 1666464484
transform 1 0 36667 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_141
timestamp 1666464484
transform 1 0 36655 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_142
timestamp 1666464484
transform 1 0 36667 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_143
timestamp 1666464484
transform 1 0 36737 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_144
timestamp 1666464484
transform 1 0 35419 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_145
timestamp 1666464484
transform 1 0 35407 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_146
timestamp 1666464484
transform 1 0 35419 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_147
timestamp 1666464484
transform 1 0 35489 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_148
timestamp 1666464484
transform 1 0 34171 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_149
timestamp 1666464484
transform 1 0 34159 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_150
timestamp 1666464484
transform 1 0 34171 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_151
timestamp 1666464484
transform 1 0 34241 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_152
timestamp 1666464484
transform 1 0 32923 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_153
timestamp 1666464484
transform 1 0 32911 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_154
timestamp 1666464484
transform 1 0 32923 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_155
timestamp 1666464484
transform 1 0 32993 0 1 2010
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_156
timestamp 1666464484
transform 1 0 31675 0 1 398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_157
timestamp 1666464484
transform 1 0 31663 0 1 1236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_158
timestamp 1666464484
transform 1 0 31675 0 1 76
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_159
timestamp 1666464484
transform 1 0 31745 0 1 2010
box 0 0 1 1
<< labels >>
rlabel metal3 s 21744 1993 21842 2091 4 gnd
port 1 nsew
rlabel metal3 s 26736 1993 26834 2091 4 gnd
port 1 nsew
rlabel metal3 s 32976 1993 33074 2091 4 gnd
port 1 nsew
rlabel metal3 s 24240 1993 24338 2091 4 gnd
port 1 nsew
rlabel metal3 s 29232 1993 29330 2091 4 gnd
port 1 nsew
rlabel metal3 s 40464 1993 40562 2091 4 gnd
port 1 nsew
rlabel metal3 s 35472 1993 35570 2091 4 gnd
port 1 nsew
rlabel metal3 s 25488 1993 25586 2091 4 gnd
port 1 nsew
rlabel metal3 s 34224 1993 34322 2091 4 gnd
port 1 nsew
rlabel metal3 s 37968 1993 38066 2091 4 gnd
port 1 nsew
rlabel metal3 s 30480 1993 30578 2091 4 gnd
port 1 nsew
rlabel metal3 s 31728 1993 31826 2091 4 gnd
port 1 nsew
rlabel metal3 s 39216 1993 39314 2091 4 gnd
port 1 nsew
rlabel metal3 s 36720 1993 36818 2091 4 gnd
port 1 nsew
rlabel metal3 s 27984 1993 28082 2091 4 gnd
port 1 nsew
rlabel metal3 s 22992 1993 23090 2091 4 gnd
port 1 nsew
rlabel metal3 s 39146 381 39244 479 4 vdd
port 2 nsew
rlabel metal3 s 22922 381 23020 479 4 vdd
port 2 nsew
rlabel metal3 s 32894 1219 32992 1317 4 vdd
port 2 nsew
rlabel metal3 s 34142 1219 34240 1317 4 vdd
port 2 nsew
rlabel metal3 s 35402 381 35500 479 4 vdd
port 2 nsew
rlabel metal3 s 37898 381 37996 479 4 vdd
port 2 nsew
rlabel metal3 s 25418 381 25516 479 4 vdd
port 2 nsew
rlabel metal3 s 26654 1219 26752 1317 4 vdd
port 2 nsew
rlabel metal3 s 27914 381 28012 479 4 vdd
port 2 nsew
rlabel metal3 s 36638 1219 36736 1317 4 vdd
port 2 nsew
rlabel metal3 s 40394 381 40492 479 4 vdd
port 2 nsew
rlabel metal3 s 24170 381 24268 479 4 vdd
port 2 nsew
rlabel metal3 s 22910 1219 23008 1317 4 vdd
port 2 nsew
rlabel metal3 s 36650 381 36748 479 4 vdd
port 2 nsew
rlabel metal3 s 25406 1219 25504 1317 4 vdd
port 2 nsew
rlabel metal3 s 32906 381 33004 479 4 vdd
port 2 nsew
rlabel metal3 s 35390 1219 35488 1317 4 vdd
port 2 nsew
rlabel metal3 s 29162 381 29260 479 4 vdd
port 2 nsew
rlabel metal3 s 21662 1219 21760 1317 4 vdd
port 2 nsew
rlabel metal3 s 27902 1219 28000 1317 4 vdd
port 2 nsew
rlabel metal3 s 31646 1219 31744 1317 4 vdd
port 2 nsew
rlabel metal3 s 24158 1219 24256 1317 4 vdd
port 2 nsew
rlabel metal3 s 30398 1219 30496 1317 4 vdd
port 2 nsew
rlabel metal3 s 37886 1219 37984 1317 4 vdd
port 2 nsew
rlabel metal3 s 26666 381 26764 479 4 vdd
port 2 nsew
rlabel metal3 s 30410 381 30508 479 4 vdd
port 2 nsew
rlabel metal3 s 31658 381 31756 479 4 vdd
port 2 nsew
rlabel metal3 s 34154 381 34252 479 4 vdd
port 2 nsew
rlabel metal3 s 40382 1219 40480 1317 4 vdd
port 2 nsew
rlabel metal3 s 21674 381 21772 479 4 vdd
port 2 nsew
rlabel metal3 s 29150 1219 29248 1317 4 vdd
port 2 nsew
rlabel metal3 s 39134 1219 39232 1317 4 vdd
port 2 nsew
rlabel metal3 s 8016 1993 8114 2091 4 gnd
port 1 nsew
rlabel metal3 s 6686 1219 6784 1317 4 vdd
port 2 nsew
rlabel metal3 s 2954 381 3052 479 4 vdd
port 2 nsew
rlabel metal3 s 11678 1219 11776 1317 4 vdd
port 2 nsew
rlabel metal3 s 14186 381 14284 479 4 vdd
port 2 nsew
rlabel metal3 s 16682 381 16780 479 4 vdd
port 2 nsew
rlabel metal3 s 9264 1993 9362 2091 4 gnd
port 1 nsew
rlabel metal3 s 15504 1993 15602 2091 4 gnd
port 1 nsew
rlabel metal3 s 18000 1993 18098 2091 4 gnd
port 1 nsew
rlabel metal3 s 4272 1993 4370 2091 4 gnd
port 1 nsew
rlabel metal3 s 13008 1993 13106 2091 4 gnd
port 1 nsew
rlabel metal3 s 1776 1993 1874 2091 4 gnd
port 1 nsew
rlabel metal3 s 6768 1993 6866 2091 4 gnd
port 1 nsew
rlabel metal3 s 20496 1993 20594 2091 4 gnd
port 1 nsew
rlabel metal3 s 19248 1993 19346 2091 4 gnd
port 1 nsew
rlabel metal3 s 11760 1993 11858 2091 4 gnd
port 1 nsew
rlabel metal3 s 14174 1219 14272 1317 4 vdd
port 2 nsew
rlabel metal3 s 2942 1219 3040 1317 4 vdd
port 2 nsew
rlabel metal3 s 12926 1219 13024 1317 4 vdd
port 2 nsew
rlabel metal3 s 17930 381 18028 479 4 vdd
port 2 nsew
rlabel metal3 s 19178 381 19276 479 4 vdd
port 2 nsew
rlabel metal3 s 15422 1219 15520 1317 4 vdd
port 2 nsew
rlabel metal3 s 3024 1993 3122 2091 4 gnd
port 1 nsew
rlabel metal3 s 1706 381 1804 479 4 vdd
port 2 nsew
rlabel metal3 s 5450 381 5548 479 4 vdd
port 2 nsew
rlabel metal3 s 19166 1219 19264 1317 4 vdd
port 2 nsew
rlabel metal3 s 4190 1219 4288 1317 4 vdd
port 2 nsew
rlabel metal3 s 14256 1993 14354 2091 4 gnd
port 1 nsew
rlabel metal3 s 16670 1219 16768 1317 4 vdd
port 2 nsew
rlabel metal3 s 20414 1219 20512 1317 4 vdd
port 2 nsew
rlabel metal3 s 12938 381 13036 479 4 vdd
port 2 nsew
rlabel metal3 s 20426 381 20524 479 4 vdd
port 2 nsew
rlabel metal3 s 10512 1993 10610 2091 4 gnd
port 1 nsew
rlabel metal3 s 10442 381 10540 479 4 vdd
port 2 nsew
rlabel metal3 s 7934 1219 8032 1317 4 vdd
port 2 nsew
rlabel metal3 s 4202 381 4300 479 4 vdd
port 2 nsew
rlabel metal3 s 5520 1993 5618 2091 4 gnd
port 1 nsew
rlabel metal3 s 17918 1219 18016 1317 4 vdd
port 2 nsew
rlabel metal3 s 16752 1993 16850 2091 4 gnd
port 1 nsew
rlabel metal3 s 11690 381 11788 479 4 vdd
port 2 nsew
rlabel metal3 s 5438 1219 5536 1317 4 vdd
port 2 nsew
rlabel metal3 s 6698 381 6796 479 4 vdd
port 2 nsew
rlabel metal3 s 7946 381 8044 479 4 vdd
port 2 nsew
rlabel metal3 s 9194 381 9292 479 4 vdd
port 2 nsew
rlabel metal3 s 9182 1219 9280 1317 4 vdd
port 2 nsew
rlabel metal3 s 1694 1219 1792 1317 4 vdd
port 2 nsew
rlabel metal3 s 10430 1219 10528 1317 4 vdd
port 2 nsew
rlabel metal3 s 15434 381 15532 479 4 vdd
port 2 nsew
rlabel metal3 s 0 2164 40562 2224 4 en
port 3 nsew
rlabel metal3 s 15434 59 15532 157 4 gnd
port 1 nsew
rlabel metal3 s 20426 59 20524 157 4 gnd
port 1 nsew
rlabel metal3 s 19178 59 19276 157 4 gnd
port 1 nsew
rlabel metal3 s 16682 59 16780 157 4 gnd
port 1 nsew
rlabel metal3 s 4202 59 4300 157 4 gnd
port 1 nsew
rlabel metal3 s 17930 59 18028 157 4 gnd
port 1 nsew
rlabel metal3 s 5450 59 5548 157 4 gnd
port 1 nsew
rlabel metal3 s 1706 59 1804 157 4 gnd
port 1 nsew
rlabel metal3 s 12938 59 13036 157 4 gnd
port 1 nsew
rlabel metal3 s 9194 59 9292 157 4 gnd
port 1 nsew
rlabel metal3 s 10442 59 10540 157 4 gnd
port 1 nsew
rlabel metal3 s 6698 59 6796 157 4 gnd
port 1 nsew
rlabel metal3 s 11690 59 11788 157 4 gnd
port 1 nsew
rlabel metal3 s 14186 59 14284 157 4 gnd
port 1 nsew
rlabel metal3 s 2954 59 3052 157 4 gnd
port 1 nsew
rlabel metal3 s 7946 59 8044 157 4 gnd
port 1 nsew
rlabel metal3 s 32906 59 33004 157 4 gnd
port 1 nsew
rlabel metal3 s 25418 59 25516 157 4 gnd
port 1 nsew
rlabel metal3 s 37898 59 37996 157 4 gnd
port 1 nsew
rlabel metal3 s 31658 59 31756 157 4 gnd
port 1 nsew
rlabel metal3 s 27914 59 28012 157 4 gnd
port 1 nsew
rlabel metal3 s 39146 59 39244 157 4 gnd
port 1 nsew
rlabel metal3 s 36650 59 36748 157 4 gnd
port 1 nsew
rlabel metal3 s 26666 59 26764 157 4 gnd
port 1 nsew
rlabel metal3 s 21674 59 21772 157 4 gnd
port 1 nsew
rlabel metal3 s 40394 59 40492 157 4 gnd
port 1 nsew
rlabel metal3 s 35402 59 35500 157 4 gnd
port 1 nsew
rlabel metal3 s 22922 59 23020 157 4 gnd
port 1 nsew
rlabel metal3 s 29162 59 29260 157 4 gnd
port 1 nsew
rlabel metal3 s 30410 59 30508 157 4 gnd
port 1 nsew
rlabel metal3 s 24170 59 24268 157 4 gnd
port 1 nsew
rlabel metal3 s 34154 59 34252 157 4 gnd
port 1 nsew
rlabel metal1 s 1570 1130 1604 2256 4 bl_0
port 4 nsew
rlabel metal1 s 1646 1142 1674 2256 4 br_0
port 5 nsew
rlabel metal1 s 1478 0 1524 254 4 data_0
port 6 nsew
rlabel metal1 s 2818 1130 2852 2256 4 bl_1
port 7 nsew
rlabel metal1 s 2894 1142 2922 2256 4 br_1
port 8 nsew
rlabel metal1 s 2726 0 2772 254 4 data_1
port 9 nsew
rlabel metal1 s 4066 1130 4100 2256 4 bl_2
port 10 nsew
rlabel metal1 s 4142 1142 4170 2256 4 br_2
port 11 nsew
rlabel metal1 s 3974 0 4020 254 4 data_2
port 12 nsew
rlabel metal1 s 5314 1130 5348 2256 4 bl_3
port 13 nsew
rlabel metal1 s 5390 1142 5418 2256 4 br_3
port 14 nsew
rlabel metal1 s 5222 0 5268 254 4 data_3
port 15 nsew
rlabel metal1 s 6562 1130 6596 2256 4 bl_4
port 16 nsew
rlabel metal1 s 6638 1142 6666 2256 4 br_4
port 17 nsew
rlabel metal1 s 6470 0 6516 254 4 data_4
port 18 nsew
rlabel metal1 s 7810 1130 7844 2256 4 bl_5
port 19 nsew
rlabel metal1 s 7886 1142 7914 2256 4 br_5
port 20 nsew
rlabel metal1 s 7718 0 7764 254 4 data_5
port 21 nsew
rlabel metal1 s 9058 1130 9092 2256 4 bl_6
port 22 nsew
rlabel metal1 s 9134 1142 9162 2256 4 br_6
port 23 nsew
rlabel metal1 s 8966 0 9012 254 4 data_6
port 24 nsew
rlabel metal1 s 10306 1130 10340 2256 4 bl_7
port 25 nsew
rlabel metal1 s 10382 1142 10410 2256 4 br_7
port 26 nsew
rlabel metal1 s 10214 0 10260 254 4 data_7
port 27 nsew
rlabel metal1 s 11554 1130 11588 2256 4 bl_8
port 28 nsew
rlabel metal1 s 11630 1142 11658 2256 4 br_8
port 29 nsew
rlabel metal1 s 11462 0 11508 254 4 data_8
port 30 nsew
rlabel metal1 s 12802 1130 12836 2256 4 bl_9
port 31 nsew
rlabel metal1 s 12878 1142 12906 2256 4 br_9
port 32 nsew
rlabel metal1 s 12710 0 12756 254 4 data_9
port 33 nsew
rlabel metal1 s 14050 1130 14084 2256 4 bl_10
port 34 nsew
rlabel metal1 s 14126 1142 14154 2256 4 br_10
port 35 nsew
rlabel metal1 s 13958 0 14004 254 4 data_10
port 36 nsew
rlabel metal1 s 15298 1130 15332 2256 4 bl_11
port 37 nsew
rlabel metal1 s 15374 1142 15402 2256 4 br_11
port 38 nsew
rlabel metal1 s 15206 0 15252 254 4 data_11
port 39 nsew
rlabel metal1 s 16546 1130 16580 2256 4 bl_12
port 40 nsew
rlabel metal1 s 16622 1142 16650 2256 4 br_12
port 41 nsew
rlabel metal1 s 16454 0 16500 254 4 data_12
port 42 nsew
rlabel metal1 s 17794 1130 17828 2256 4 bl_13
port 43 nsew
rlabel metal1 s 17870 1142 17898 2256 4 br_13
port 44 nsew
rlabel metal1 s 17702 0 17748 254 4 data_13
port 45 nsew
rlabel metal1 s 19042 1130 19076 2256 4 bl_14
port 46 nsew
rlabel metal1 s 19118 1142 19146 2256 4 br_14
port 47 nsew
rlabel metal1 s 18950 0 18996 254 4 data_14
port 48 nsew
rlabel metal1 s 20290 1130 20324 2256 4 bl_15
port 49 nsew
rlabel metal1 s 20366 1142 20394 2256 4 br_15
port 50 nsew
rlabel metal1 s 20198 0 20244 254 4 data_15
port 51 nsew
rlabel metal1 s 21538 1130 21572 2256 4 bl_16
port 52 nsew
rlabel metal1 s 21614 1142 21642 2256 4 br_16
port 53 nsew
rlabel metal1 s 21446 0 21492 254 4 data_16
port 54 nsew
rlabel metal1 s 22786 1130 22820 2256 4 bl_17
port 55 nsew
rlabel metal1 s 22862 1142 22890 2256 4 br_17
port 56 nsew
rlabel metal1 s 22694 0 22740 254 4 data_17
port 57 nsew
rlabel metal1 s 24034 1130 24068 2256 4 bl_18
port 58 nsew
rlabel metal1 s 24110 1142 24138 2256 4 br_18
port 59 nsew
rlabel metal1 s 23942 0 23988 254 4 data_18
port 60 nsew
rlabel metal1 s 25282 1130 25316 2256 4 bl_19
port 61 nsew
rlabel metal1 s 25358 1142 25386 2256 4 br_19
port 62 nsew
rlabel metal1 s 25190 0 25236 254 4 data_19
port 63 nsew
rlabel metal1 s 26530 1130 26564 2256 4 bl_20
port 64 nsew
rlabel metal1 s 26606 1142 26634 2256 4 br_20
port 65 nsew
rlabel metal1 s 26438 0 26484 254 4 data_20
port 66 nsew
rlabel metal1 s 27778 1130 27812 2256 4 bl_21
port 67 nsew
rlabel metal1 s 27854 1142 27882 2256 4 br_21
port 68 nsew
rlabel metal1 s 27686 0 27732 254 4 data_21
port 69 nsew
rlabel metal1 s 29026 1130 29060 2256 4 bl_22
port 70 nsew
rlabel metal1 s 29102 1142 29130 2256 4 br_22
port 71 nsew
rlabel metal1 s 28934 0 28980 254 4 data_22
port 72 nsew
rlabel metal1 s 30274 1130 30308 2256 4 bl_23
port 73 nsew
rlabel metal1 s 30350 1142 30378 2256 4 br_23
port 74 nsew
rlabel metal1 s 30182 0 30228 254 4 data_23
port 75 nsew
rlabel metal1 s 31522 1130 31556 2256 4 bl_24
port 76 nsew
rlabel metal1 s 31598 1142 31626 2256 4 br_24
port 77 nsew
rlabel metal1 s 31430 0 31476 254 4 data_24
port 78 nsew
rlabel metal1 s 32770 1130 32804 2256 4 bl_25
port 79 nsew
rlabel metal1 s 32846 1142 32874 2256 4 br_25
port 80 nsew
rlabel metal1 s 32678 0 32724 254 4 data_25
port 81 nsew
rlabel metal1 s 34018 1130 34052 2256 4 bl_26
port 82 nsew
rlabel metal1 s 34094 1142 34122 2256 4 br_26
port 83 nsew
rlabel metal1 s 33926 0 33972 254 4 data_26
port 84 nsew
rlabel metal1 s 35266 1130 35300 2256 4 bl_27
port 85 nsew
rlabel metal1 s 35342 1142 35370 2256 4 br_27
port 86 nsew
rlabel metal1 s 35174 0 35220 254 4 data_27
port 87 nsew
rlabel metal1 s 36514 1130 36548 2256 4 bl_28
port 88 nsew
rlabel metal1 s 36590 1142 36618 2256 4 br_28
port 89 nsew
rlabel metal1 s 36422 0 36468 254 4 data_28
port 90 nsew
rlabel metal1 s 37762 1130 37796 2256 4 bl_29
port 91 nsew
rlabel metal1 s 37838 1142 37866 2256 4 br_29
port 92 nsew
rlabel metal1 s 37670 0 37716 254 4 data_29
port 93 nsew
rlabel metal1 s 39010 1130 39044 2256 4 bl_30
port 94 nsew
rlabel metal1 s 39086 1142 39114 2256 4 br_30
port 95 nsew
rlabel metal1 s 38918 0 38964 254 4 data_30
port 96 nsew
rlabel metal1 s 40258 1130 40292 2256 4 bl_31
port 97 nsew
rlabel metal1 s 40334 1142 40362 2256 4 br_31
port 98 nsew
rlabel metal1 s 40166 0 40212 254 4 data_31
port 99 nsew
<< properties >>
string FIXED_BBOX 0 0 40562 2256
string GDS_END 1271198
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 1195690
<< end >>
