magic
tech sky130B
magscale 1 2
timestamp 1672577215
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 170306 700680 170312 700732
rect 170364 700720 170370 700732
rect 178310 700720 178316 700732
rect 170364 700692 178316 700720
rect 170364 700680 170370 700692
rect 178310 700680 178316 700692
rect 178368 700680 178374 700732
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 178402 700652 178408 700664
rect 154172 700624 178408 700652
rect 154172 700612 154178 700624
rect 178402 700612 178408 700624
rect 178460 700612 178466 700664
rect 137830 700544 137836 700596
rect 137888 700584 137894 700596
rect 178034 700584 178040 700596
rect 137888 700556 178040 700584
rect 137888 700544 137894 700556
rect 178034 700544 178040 700556
rect 178092 700544 178098 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 178218 700516 178224 700528
rect 105504 700488 178224 700516
rect 105504 700476 105510 700488
rect 178218 700476 178224 700488
rect 178276 700476 178282 700528
rect 392578 700476 392584 700528
rect 392636 700516 392642 700528
rect 429838 700516 429844 700528
rect 392636 700488 429844 700516
rect 392636 700476 392642 700488
rect 429838 700476 429844 700488
rect 429896 700476 429902 700528
rect 177390 700408 177396 700460
rect 177448 700448 177454 700460
rect 283834 700448 283840 700460
rect 177448 700420 283840 700448
rect 177448 700408 177454 700420
rect 283834 700408 283840 700420
rect 283892 700408 283898 700460
rect 366358 700408 366364 700460
rect 366416 700448 366422 700460
rect 413646 700448 413652 700460
rect 366416 700420 413652 700448
rect 366416 700408 366422 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 178126 700380 178132 700392
rect 73028 700352 178132 700380
rect 73028 700340 73034 700352
rect 178126 700340 178132 700352
rect 178184 700340 178190 700392
rect 186958 700340 186964 700392
rect 187016 700380 187022 700392
rect 218974 700380 218980 700392
rect 187016 700352 218980 700380
rect 187016 700340 187022 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 360838 700340 360844 700392
rect 360896 700380 360902 700392
rect 462314 700380 462320 700392
rect 360896 700352 462320 700380
rect 360896 700340 360902 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 176654 700312 176660 700324
rect 89220 700284 176660 700312
rect 89220 700272 89226 700284
rect 176654 700272 176660 700284
rect 176712 700272 176718 700324
rect 177298 700272 177304 700324
rect 177356 700312 177362 700324
rect 348786 700312 348792 700324
rect 177356 700284 348792 700312
rect 177356 700272 177362 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 363598 700272 363604 700324
rect 363656 700312 363662 700324
rect 478506 700312 478512 700324
rect 363656 700284 478512 700312
rect 363656 700272 363662 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 26878 699700 26884 699712
rect 24360 699672 26884 699700
rect 24360 699660 24366 699672
rect 26878 699660 26884 699672
rect 26936 699660 26942 699712
rect 192478 696940 192484 696992
rect 192536 696980 192542 696992
rect 580166 696980 580172 696992
rect 192536 696952 580172 696980
rect 192536 696940 192542 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 170858 685856 170864 685908
rect 170916 685896 170922 685908
rect 192570 685896 192576 685908
rect 170916 685868 192576 685896
rect 170916 685856 170922 685868
rect 192570 685856 192576 685868
rect 192628 685856 192634 685908
rect 350994 685856 351000 685908
rect 351052 685896 351058 685908
rect 378778 685896 378784 685908
rect 351052 685868 378784 685896
rect 351052 685856 351058 685868
rect 378778 685856 378784 685868
rect 378836 685856 378842 685908
rect 530946 685856 530952 685908
rect 531004 685896 531010 685908
rect 536834 685896 536840 685908
rect 531004 685868 536840 685896
rect 531004 685856 531010 685868
rect 536834 685856 536840 685868
rect 536892 685856 536898 685908
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 18598 683176 18604 683188
rect 3476 683148 18604 683176
rect 3476 683136 3482 683148
rect 18598 683136 18604 683148
rect 18656 683136 18662 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 18690 670732 18696 670744
rect 3568 670704 18696 670732
rect 3568 670692 3574 670704
rect 18690 670692 18696 670704
rect 18748 670692 18754 670744
rect 538858 670692 538864 670744
rect 538916 670732 538922 670744
rect 580166 670732 580172 670744
rect 538916 670704 580172 670732
rect 538916 670692 538922 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 31018 656928 31024 656940
rect 3476 656900 31024 656928
rect 3476 656888 3482 656900
rect 31018 656888 31024 656900
rect 31076 656888 31082 656940
rect 537478 643084 537484 643136
rect 537536 643124 537542 643136
rect 580166 643124 580172 643136
rect 537536 643096 580172 643124
rect 537536 643084 537542 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 25498 618304 25504 618316
rect 3200 618276 25504 618304
rect 3200 618264 3206 618276
rect 25498 618264 25504 618276
rect 25556 618264 25562 618316
rect 538950 616836 538956 616888
rect 539008 616876 539014 616888
rect 580166 616876 580172 616888
rect 539008 616848 580172 616876
rect 539008 616836 539014 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 192570 607860 192576 607912
rect 192628 607900 192634 607912
rect 213914 607900 213920 607912
rect 192628 607872 213920 607900
rect 192628 607860 192634 607872
rect 213914 607860 213920 607872
rect 213972 607860 213978 607912
rect 378778 607860 378784 607912
rect 378836 607900 378842 607912
rect 394694 607900 394700 607912
rect 378836 607872 394700 607900
rect 378836 607860 378842 607872
rect 394694 607860 394700 607872
rect 394752 607860 394758 607912
rect 213914 607316 213920 607368
rect 213972 607356 213978 607368
rect 216674 607356 216680 607368
rect 213972 607328 216680 607356
rect 213972 607316 213978 607328
rect 216674 607316 216680 607328
rect 216732 607316 216738 607368
rect 394694 607180 394700 607232
rect 394752 607220 394758 607232
rect 397178 607220 397184 607232
rect 394752 607192 397184 607220
rect 394752 607180 394758 607192
rect 397178 607180 397184 607192
rect 397236 607180 397242 607232
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 11698 605860 11704 605872
rect 3292 605832 11704 605860
rect 3292 605820 3298 605832
rect 11698 605820 11704 605832
rect 11756 605820 11762 605872
rect 66806 597456 66812 597508
rect 66864 597496 66870 597508
rect 84194 597496 84200 597508
rect 66864 597468 84200 597496
rect 66864 597456 66870 597468
rect 84194 597456 84200 597468
rect 84252 597456 84258 597508
rect 397730 597456 397736 597508
rect 397788 597496 397794 597508
rect 436002 597496 436008 597508
rect 397788 597468 436008 597496
rect 397788 597456 397794 597468
rect 436002 597456 436008 597468
rect 436060 597456 436066 597508
rect 74902 597388 74908 597440
rect 74960 597428 74966 597440
rect 92474 597428 92480 597440
rect 74960 597400 92480 597428
rect 74960 597388 74966 597400
rect 92474 597388 92480 597400
rect 92532 597388 92538 597440
rect 399478 597388 399484 597440
rect 399536 597428 399542 597440
rect 434622 597428 434628 597440
rect 399536 597400 434628 597428
rect 399536 597388 399542 597400
rect 434622 597388 434628 597400
rect 434680 597388 434686 597440
rect 68738 597320 68744 597372
rect 68796 597360 68802 597372
rect 85574 597360 85580 597372
rect 68796 597332 85580 597360
rect 68796 597320 68802 597332
rect 85574 597320 85580 597332
rect 85632 597320 85638 597372
rect 397822 597320 397828 597372
rect 397880 597360 397886 597372
rect 437106 597360 437112 597372
rect 397880 597332 437112 597360
rect 397880 597320 397886 597332
rect 437106 597320 437112 597332
rect 437164 597320 437170 597372
rect 66162 597252 66168 597304
rect 66220 597292 66226 597304
rect 82814 597292 82820 597304
rect 66220 597264 82820 597292
rect 66220 597252 66226 597264
rect 82814 597252 82820 597264
rect 82872 597252 82878 597304
rect 395338 597252 395344 597304
rect 395396 597292 395402 597304
rect 434714 597292 434720 597304
rect 395396 597264 434720 597292
rect 395396 597252 395402 597264
rect 434714 597252 434720 597264
rect 434772 597252 434778 597304
rect 39206 597184 39212 597236
rect 39264 597224 39270 597236
rect 74902 597224 74908 597236
rect 39264 597196 74908 597224
rect 39264 597184 39270 597196
rect 74902 597184 74908 597196
rect 74960 597184 74966 597236
rect 77110 597184 77116 597236
rect 77168 597224 77174 597236
rect 95234 597224 95240 597236
rect 77168 597196 95240 597224
rect 77168 597184 77174 597196
rect 95234 597184 95240 597196
rect 95292 597184 95298 597236
rect 256694 597184 256700 597236
rect 256752 597224 256758 597236
rect 274634 597224 274640 597236
rect 256752 597196 274640 597224
rect 256752 597184 256758 597196
rect 274634 597184 274640 597196
rect 274692 597184 274698 597236
rect 426526 597184 426532 597236
rect 426584 597224 426590 597236
rect 444374 597224 444380 597236
rect 426584 597196 444380 597224
rect 426584 597184 426590 597196
rect 444374 597184 444380 597196
rect 444432 597184 444438 597236
rect 68830 597116 68836 597168
rect 68888 597156 68894 597168
rect 86954 597156 86960 597168
rect 68888 597128 86960 597156
rect 68888 597116 68894 597128
rect 86954 597116 86960 597128
rect 87012 597116 87018 597168
rect 214742 597116 214748 597168
rect 214800 597156 214806 597168
rect 258074 597156 258080 597168
rect 214800 597128 258080 597156
rect 214800 597116 214806 597128
rect 258074 597116 258080 597128
rect 258132 597156 258138 597168
rect 276014 597156 276020 597168
rect 258132 597128 276020 597156
rect 258132 597116 258138 597128
rect 276014 597116 276020 597128
rect 276072 597116 276078 597168
rect 425606 597116 425612 597168
rect 425664 597156 425670 597168
rect 443638 597156 443644 597168
rect 425664 597128 443644 597156
rect 425664 597116 425670 597128
rect 443638 597116 443644 597128
rect 443696 597116 443702 597168
rect 36906 597048 36912 597100
rect 36964 597088 36970 597100
rect 78030 597088 78036 597100
rect 36964 597060 78036 597088
rect 36964 597048 36970 597060
rect 78030 597048 78036 597060
rect 78088 597088 78094 597100
rect 96614 597088 96620 597100
rect 78088 597060 96620 597088
rect 78088 597048 78094 597060
rect 96614 597048 96620 597060
rect 96672 597048 96678 597100
rect 139302 597048 139308 597100
rect 139360 597088 139366 597100
rect 178954 597088 178960 597100
rect 139360 597060 178960 597088
rect 139360 597048 139366 597060
rect 178954 597048 178960 597060
rect 179012 597048 179018 597100
rect 243078 597048 243084 597100
rect 243136 597088 243142 597100
rect 260834 597088 260840 597100
rect 243136 597060 260840 597088
rect 243136 597048 243142 597060
rect 260834 597048 260840 597060
rect 260892 597048 260898 597100
rect 424962 597048 424968 597100
rect 425020 597088 425026 597100
rect 441982 597088 441988 597100
rect 425020 597060 441988 597088
rect 425020 597048 425026 597060
rect 441982 597048 441988 597060
rect 442040 597048 442046 597100
rect 39942 596980 39948 597032
rect 40000 597020 40006 597032
rect 56594 597020 56600 597032
rect 40000 596992 56600 597020
rect 40000 596980 40006 596992
rect 56594 596980 56600 596992
rect 56652 596980 56658 597032
rect 69750 596980 69756 597032
rect 69808 597020 69814 597032
rect 88334 597020 88340 597032
rect 69808 596992 88340 597020
rect 69808 596980 69814 596992
rect 88334 596980 88340 596992
rect 88392 596980 88398 597032
rect 126882 596980 126888 597032
rect 126940 597020 126946 597032
rect 177942 597020 177948 597032
rect 126940 596992 177948 597020
rect 126940 596980 126946 596992
rect 177942 596980 177948 596992
rect 178000 596980 178006 597032
rect 219710 596980 219716 597032
rect 219768 597020 219774 597032
rect 235994 597020 236000 597032
rect 219768 596992 236000 597020
rect 219768 596980 219774 596992
rect 235994 596980 236000 596992
rect 236052 596980 236058 597032
rect 244274 596980 244280 597032
rect 244332 597020 244338 597032
rect 262214 597020 262220 597032
rect 244332 596992 262220 597020
rect 244332 596980 244338 596992
rect 262214 596980 262220 596992
rect 262272 596980 262278 597032
rect 399662 596980 399668 597032
rect 399720 597020 399726 597032
rect 416774 597020 416780 597032
rect 399720 596992 416780 597020
rect 399720 596980 399726 596992
rect 416774 596980 416780 596992
rect 416832 596980 416838 597032
rect 434622 596980 434628 597032
rect 434680 597020 434686 597032
rect 452654 597020 452660 597032
rect 434680 596992 452660 597020
rect 434680 596980 434686 596992
rect 452654 596980 452660 596992
rect 452712 596980 452718 597032
rect 39666 596912 39672 596964
rect 39724 596952 39730 596964
rect 59354 596952 59360 596964
rect 39724 596924 59360 596952
rect 39724 596912 39730 596924
rect 59354 596912 59360 596924
rect 59412 596912 59418 596964
rect 70394 596912 70400 596964
rect 70452 596952 70458 596964
rect 71314 596952 71320 596964
rect 70452 596924 71320 596952
rect 70452 596912 70458 596924
rect 71314 596912 71320 596924
rect 71372 596952 71378 596964
rect 89714 596952 89720 596964
rect 71372 596924 89720 596952
rect 71372 596912 71378 596924
rect 89714 596912 89720 596924
rect 89772 596912 89778 596964
rect 118602 596912 118608 596964
rect 118660 596952 118666 596964
rect 178770 596952 178776 596964
rect 118660 596924 178776 596952
rect 118660 596912 118666 596924
rect 178770 596912 178776 596924
rect 178828 596912 178834 596964
rect 218882 596912 218888 596964
rect 218940 596952 218946 596964
rect 236178 596952 236184 596964
rect 218940 596924 236184 596952
rect 218940 596912 218946 596924
rect 236178 596912 236184 596924
rect 236236 596912 236242 596964
rect 244366 596912 244372 596964
rect 244424 596952 244430 596964
rect 245470 596952 245476 596964
rect 244424 596924 245476 596952
rect 244424 596912 244430 596924
rect 245470 596912 245476 596924
rect 245528 596952 245534 596964
rect 263686 596952 263692 596964
rect 245528 596924 263692 596952
rect 245528 596912 245534 596924
rect 263686 596912 263692 596924
rect 263744 596912 263750 596964
rect 399938 596912 399944 596964
rect 399996 596952 400002 596964
rect 419534 596952 419540 596964
rect 399996 596924 419540 596952
rect 399996 596912 400002 596924
rect 419534 596912 419540 596924
rect 419592 596912 419598 596964
rect 436002 596912 436008 596964
rect 436060 596952 436066 596964
rect 454034 596952 454040 596964
rect 436060 596924 454040 596952
rect 436060 596912 436066 596924
rect 454034 596912 454040 596924
rect 454092 596912 454098 596964
rect 39482 596844 39488 596896
rect 39540 596884 39546 596896
rect 63218 596884 63224 596896
rect 39540 596856 63224 596884
rect 39540 596844 39546 596856
rect 63218 596844 63224 596856
rect 63276 596884 63282 596896
rect 81434 596884 81440 596896
rect 63276 596856 81440 596884
rect 63276 596844 63282 596856
rect 81434 596844 81440 596856
rect 81492 596844 81498 596896
rect 121362 596844 121368 596896
rect 121420 596884 121426 596896
rect 182818 596884 182824 596896
rect 121420 596856 182824 596884
rect 121420 596844 121426 596856
rect 182818 596844 182824 596856
rect 182876 596844 182882 596896
rect 219066 596844 219072 596896
rect 219124 596884 219130 596896
rect 237374 596884 237380 596896
rect 219124 596856 237380 596884
rect 219124 596844 219130 596856
rect 237374 596844 237380 596856
rect 237432 596844 237438 596896
rect 253934 596844 253940 596896
rect 253992 596884 253998 596896
rect 254578 596884 254584 596896
rect 253992 596856 254584 596884
rect 253992 596844 253998 596856
rect 254578 596844 254584 596856
rect 254636 596884 254642 596896
rect 273254 596884 273260 596896
rect 254636 596856 273260 596884
rect 254636 596844 254642 596856
rect 273254 596844 273260 596856
rect 273312 596844 273318 596896
rect 326982 596844 326988 596896
rect 327040 596884 327046 596896
rect 358998 596884 359004 596896
rect 327040 596856 359004 596884
rect 327040 596844 327046 596856
rect 358998 596844 359004 596856
rect 359056 596844 359062 596896
rect 398282 596844 398288 596896
rect 398340 596884 398346 596896
rect 418154 596884 418160 596896
rect 398340 596856 418160 596884
rect 398340 596844 398346 596856
rect 418154 596844 418160 596856
rect 418212 596844 418218 596896
rect 437106 596844 437112 596896
rect 437164 596884 437170 596896
rect 455414 596884 455420 596896
rect 437164 596856 455420 596884
rect 437164 596844 437170 596856
rect 455414 596844 455420 596856
rect 455472 596844 455478 596896
rect 39758 596776 39764 596828
rect 39816 596816 39822 596828
rect 64230 596816 64236 596828
rect 39816 596788 64236 596816
rect 39816 596776 39822 596788
rect 64230 596776 64236 596788
rect 64288 596816 64294 596828
rect 82814 596816 82820 596828
rect 64288 596788 82820 596816
rect 64288 596776 64294 596788
rect 82814 596776 82820 596788
rect 82872 596776 82878 596828
rect 117222 596776 117228 596828
rect 117280 596816 117286 596828
rect 178862 596816 178868 596828
rect 117280 596788 178868 596816
rect 117280 596776 117286 596788
rect 178862 596776 178868 596788
rect 178920 596776 178926 596828
rect 219250 596776 219256 596828
rect 219308 596816 219314 596828
rect 238754 596816 238760 596828
rect 219308 596788 238760 596816
rect 219308 596776 219314 596788
rect 238754 596776 238760 596788
rect 238812 596776 238818 596828
rect 245654 596776 245660 596828
rect 245712 596816 245718 596828
rect 246482 596816 246488 596828
rect 245712 596788 246488 596816
rect 245712 596776 245718 596788
rect 246482 596776 246488 596788
rect 246540 596816 246546 596828
rect 265066 596816 265072 596828
rect 246540 596788 265072 596816
rect 246540 596776 246546 596788
rect 265066 596776 265072 596788
rect 265124 596776 265130 596828
rect 324222 596776 324228 596828
rect 324280 596816 324286 596828
rect 357894 596816 357900 596828
rect 324280 596788 357900 596816
rect 324280 596776 324286 596788
rect 357894 596776 357900 596788
rect 357952 596776 357958 596828
rect 398558 596776 398564 596828
rect 398616 596816 398622 596828
rect 419534 596816 419540 596828
rect 398616 596788 419540 596816
rect 398616 596776 398622 596788
rect 419534 596776 419540 596788
rect 419592 596776 419598 596828
rect 423122 596816 423128 596828
rect 422266 596788 423128 596816
rect 38378 596708 38384 596760
rect 38436 596748 38442 596760
rect 64874 596748 64880 596760
rect 38436 596720 64880 596748
rect 38436 596708 38442 596720
rect 64874 596708 64880 596720
rect 64932 596748 64938 596760
rect 66162 596748 66168 596760
rect 64932 596720 66168 596748
rect 64932 596708 64938 596720
rect 66162 596708 66168 596720
rect 66220 596708 66226 596760
rect 114462 596708 114468 596760
rect 114520 596748 114526 596760
rect 178678 596748 178684 596760
rect 114520 596720 178684 596748
rect 114520 596708 114526 596720
rect 178678 596708 178684 596720
rect 178736 596708 178742 596760
rect 218974 596708 218980 596760
rect 219032 596748 219038 596760
rect 240134 596748 240140 596760
rect 219032 596720 240140 596748
rect 219032 596708 219038 596720
rect 240134 596708 240140 596720
rect 240192 596708 240198 596760
rect 252094 596708 252100 596760
rect 252152 596748 252158 596760
rect 270586 596748 270592 596760
rect 252152 596720 270592 596748
rect 252152 596708 252158 596720
rect 270586 596708 270592 596720
rect 270644 596708 270650 596760
rect 321462 596708 321468 596760
rect 321520 596748 321526 596760
rect 359090 596748 359096 596760
rect 321520 596720 359096 596748
rect 321520 596708 321526 596720
rect 359090 596708 359096 596720
rect 359148 596708 359154 596760
rect 398098 596708 398104 596760
rect 398156 596748 398162 596760
rect 420914 596748 420920 596760
rect 398156 596720 420920 596748
rect 398156 596708 398162 596720
rect 420914 596708 420920 596720
rect 420972 596708 420978 596760
rect 39390 596640 39396 596692
rect 39448 596680 39454 596692
rect 66806 596680 66812 596692
rect 39448 596652 66812 596680
rect 39448 596640 39454 596652
rect 66806 596640 66812 596652
rect 66864 596640 66870 596692
rect 111702 596640 111708 596692
rect 111760 596680 111766 596692
rect 177850 596680 177856 596692
rect 111760 596652 177856 596680
rect 111760 596640 111766 596652
rect 177850 596640 177856 596652
rect 177908 596640 177914 596692
rect 217962 596640 217968 596692
rect 218020 596680 218026 596692
rect 241514 596680 241520 596692
rect 218020 596652 241520 596680
rect 218020 596640 218026 596652
rect 241514 596640 241520 596652
rect 241572 596640 241578 596692
rect 252186 596640 252192 596692
rect 252244 596680 252250 596692
rect 269114 596680 269120 596692
rect 252244 596652 269120 596680
rect 252244 596640 252250 596652
rect 269114 596640 269120 596652
rect 269172 596640 269178 596692
rect 318702 596640 318708 596692
rect 318760 596680 318766 596692
rect 357710 596680 357716 596692
rect 318760 596652 357716 596680
rect 318760 596640 318766 596652
rect 357710 596640 357716 596652
rect 357768 596640 357774 596692
rect 399754 596640 399760 596692
rect 399812 596680 399818 596692
rect 422266 596680 422294 596788
rect 423122 596776 423128 596788
rect 423180 596816 423186 596828
rect 441614 596816 441620 596828
rect 423180 596788 441620 596816
rect 423180 596776 423186 596788
rect 441614 596776 441620 596788
rect 441672 596776 441678 596828
rect 399812 596652 422294 596680
rect 399812 596640 399818 596652
rect 39298 596572 39304 596624
rect 39356 596612 39362 596624
rect 68830 596612 68836 596624
rect 39356 596584 68836 596612
rect 39356 596572 39362 596584
rect 68830 596572 68836 596584
rect 68888 596572 68894 596624
rect 124122 596572 124128 596624
rect 124180 596612 124186 596624
rect 191098 596612 191104 596624
rect 124180 596584 191104 596612
rect 124180 596572 124186 596584
rect 191098 596572 191104 596584
rect 191156 596572 191162 596624
rect 219158 596572 219164 596624
rect 219216 596612 219222 596624
rect 243078 596612 243084 596624
rect 219216 596584 243084 596612
rect 219216 596572 219222 596584
rect 243078 596572 243084 596584
rect 243136 596572 243142 596624
rect 248414 596572 248420 596624
rect 248472 596612 248478 596624
rect 266354 596612 266360 596624
rect 248472 596584 266360 596612
rect 248472 596572 248478 596584
rect 266354 596572 266360 596584
rect 266412 596572 266418 596624
rect 314562 596572 314568 596624
rect 314620 596612 314626 596624
rect 357526 596612 357532 596624
rect 314620 596584 357532 596612
rect 314620 596572 314626 596584
rect 357526 596572 357532 596584
rect 357584 596572 357590 596624
rect 398466 596572 398472 596624
rect 398524 596612 398530 596624
rect 424962 596612 424968 596624
rect 398524 596584 424968 596612
rect 398524 596572 398530 596584
rect 424962 596572 424968 596584
rect 425020 596572 425026 596624
rect 427998 596572 428004 596624
rect 428056 596612 428062 596624
rect 447226 596612 447232 596624
rect 428056 596584 447232 596612
rect 428056 596572 428062 596584
rect 447226 596572 447232 596584
rect 447284 596572 447290 596624
rect 37642 596504 37648 596556
rect 37700 596544 37706 596556
rect 67634 596544 67640 596556
rect 37700 596516 67640 596544
rect 37700 596504 37706 596516
rect 67634 596504 67640 596516
rect 67692 596544 67698 596556
rect 68738 596544 68744 596556
rect 67692 596516 68744 596544
rect 67692 596504 67698 596516
rect 68738 596504 68744 596516
rect 68796 596504 68802 596556
rect 108942 596504 108948 596556
rect 109000 596544 109006 596556
rect 180058 596544 180064 596556
rect 109000 596516 180064 596544
rect 109000 596504 109006 596516
rect 180058 596504 180064 596516
rect 180116 596504 180122 596556
rect 218790 596504 218796 596556
rect 218848 596544 218854 596556
rect 244274 596544 244280 596556
rect 218848 596516 244280 596544
rect 218848 596504 218854 596516
rect 244274 596504 244280 596516
rect 244332 596504 244338 596556
rect 249886 596504 249892 596556
rect 249944 596544 249950 596556
rect 267918 596544 267924 596556
rect 249944 596516 267924 596544
rect 249944 596504 249950 596516
rect 267918 596504 267924 596516
rect 267976 596504 267982 596556
rect 315942 596504 315948 596556
rect 316000 596544 316006 596556
rect 359182 596544 359188 596556
rect 316000 596516 359188 596544
rect 316000 596504 316006 596516
rect 359182 596504 359188 596516
rect 359240 596504 359246 596556
rect 398374 596504 398380 596556
rect 398432 596544 398438 596556
rect 425606 596544 425612 596556
rect 398432 596516 425612 596544
rect 398432 596504 398438 596516
rect 425606 596504 425612 596516
rect 425664 596504 425670 596556
rect 426434 596504 426440 596556
rect 426492 596544 426498 596556
rect 427630 596544 427636 596556
rect 426492 596516 427636 596544
rect 426492 596504 426498 596516
rect 427630 596504 427636 596516
rect 427688 596544 427694 596556
rect 445846 596544 445852 596556
rect 427688 596516 445852 596544
rect 427688 596504 427694 596516
rect 445846 596504 445852 596516
rect 445904 596504 445910 596556
rect 37182 596436 37188 596488
rect 37240 596476 37246 596488
rect 69750 596476 69756 596488
rect 37240 596448 69756 596476
rect 37240 596436 37246 596448
rect 69750 596436 69756 596448
rect 69808 596436 69814 596488
rect 76006 596436 76012 596488
rect 76064 596476 76070 596488
rect 94038 596476 94044 596488
rect 76064 596448 94044 596476
rect 76064 596436 76070 596448
rect 94038 596436 94044 596448
rect 94096 596436 94102 596488
rect 106182 596436 106188 596488
rect 106240 596476 106246 596488
rect 177758 596476 177764 596488
rect 106240 596448 177764 596476
rect 106240 596436 106246 596448
rect 177758 596436 177764 596448
rect 177816 596436 177822 596488
rect 214834 596436 214840 596488
rect 214892 596476 214898 596488
rect 244366 596476 244372 596488
rect 214892 596448 244372 596476
rect 214892 596436 214898 596448
rect 244366 596436 244372 596448
rect 244424 596436 244430 596488
rect 247126 596436 247132 596488
rect 247184 596476 247190 596488
rect 266354 596476 266360 596488
rect 247184 596448 266360 596476
rect 247184 596436 247190 596448
rect 266354 596436 266360 596448
rect 266412 596436 266418 596488
rect 311802 596436 311808 596488
rect 311860 596476 311866 596488
rect 357618 596476 357624 596488
rect 311860 596448 357624 596476
rect 311860 596436 311866 596448
rect 357618 596436 357624 596448
rect 357676 596436 357682 596488
rect 399570 596436 399576 596488
rect 399628 596476 399634 596488
rect 426526 596476 426532 596488
rect 399628 596448 426532 596476
rect 399628 596436 399634 596448
rect 426526 596436 426532 596448
rect 426584 596436 426590 596488
rect 429194 596436 429200 596488
rect 429252 596476 429258 596488
rect 448514 596476 448520 596488
rect 429252 596448 448520 596476
rect 429252 596436 429258 596448
rect 448514 596436 448520 596448
rect 448572 596436 448578 596488
rect 37090 596368 37096 596420
rect 37148 596408 37154 596420
rect 70394 596408 70400 596420
rect 37148 596380 70400 596408
rect 37148 596368 37154 596380
rect 70394 596368 70400 596380
rect 70452 596368 70458 596420
rect 71774 596368 71780 596420
rect 71832 596408 71838 596420
rect 91094 596408 91100 596420
rect 71832 596380 91100 596408
rect 71832 596368 71838 596380
rect 91094 596368 91100 596380
rect 91152 596368 91158 596420
rect 102042 596368 102048 596420
rect 102100 596408 102106 596420
rect 177574 596408 177580 596420
rect 102100 596380 177580 596408
rect 102100 596368 102106 596380
rect 177574 596368 177580 596380
rect 177632 596368 177638 596420
rect 215110 596368 215116 596420
rect 215168 596408 215174 596420
rect 245654 596408 245660 596420
rect 215168 596380 245660 596408
rect 215168 596368 215174 596380
rect 245654 596368 245660 596380
rect 245712 596368 245718 596420
rect 253474 596368 253480 596420
rect 253532 596408 253538 596420
rect 271874 596408 271880 596420
rect 253532 596380 271880 596408
rect 253532 596368 253538 596380
rect 271874 596368 271880 596380
rect 271932 596368 271938 596420
rect 309042 596368 309048 596420
rect 309100 596408 309106 596420
rect 356606 596408 356612 596420
rect 309100 596380 356612 596408
rect 309100 596368 309106 596380
rect 356606 596368 356612 596380
rect 356664 596368 356670 596420
rect 431954 596368 431960 596420
rect 432012 596408 432018 596420
rect 449986 596408 449992 596420
rect 432012 596380 449992 596408
rect 432012 596368 432018 596380
rect 449986 596368 449992 596380
rect 450044 596368 450050 596420
rect 73154 596300 73160 596352
rect 73212 596340 73218 596352
rect 91186 596340 91192 596352
rect 73212 596312 91192 596340
rect 73212 596300 73218 596312
rect 91186 596300 91192 596312
rect 91244 596300 91250 596352
rect 99282 596300 99288 596352
rect 99340 596340 99346 596352
rect 177666 596340 177672 596352
rect 99340 596312 177672 596340
rect 99340 596300 99346 596312
rect 177666 596300 177672 596312
rect 177724 596300 177730 596352
rect 219802 596300 219808 596352
rect 219860 596340 219866 596352
rect 253934 596340 253940 596352
rect 219860 596312 253940 596340
rect 219860 596300 219866 596312
rect 253934 596300 253940 596312
rect 253992 596300 253998 596352
rect 306098 596300 306104 596352
rect 306156 596340 306162 596352
rect 357434 596340 357440 596352
rect 306156 596312 357440 596340
rect 306156 596300 306162 596312
rect 357434 596300 357440 596312
rect 357492 596300 357498 596352
rect 433426 596300 433432 596352
rect 433484 596340 433490 596352
rect 451274 596340 451280 596352
rect 433484 596312 451280 596340
rect 433484 596300 433490 596312
rect 451274 596300 451280 596312
rect 451332 596300 451338 596352
rect 37918 596232 37924 596284
rect 37976 596272 37982 596284
rect 77110 596272 77116 596284
rect 37976 596244 77116 596272
rect 37976 596232 37982 596244
rect 77110 596232 77116 596244
rect 77168 596232 77174 596284
rect 96522 596232 96528 596284
rect 96580 596272 96586 596284
rect 177482 596272 177488 596284
rect 96580 596244 177488 596272
rect 96580 596232 96586 596244
rect 177482 596232 177488 596244
rect 177540 596232 177546 596284
rect 215018 596232 215024 596284
rect 215076 596272 215082 596284
rect 256694 596272 256700 596284
rect 215076 596244 256700 596272
rect 215076 596232 215082 596244
rect 256694 596232 256700 596244
rect 256752 596232 256758 596284
rect 303522 596232 303528 596284
rect 303580 596272 303586 596284
rect 358906 596272 358912 596284
rect 303580 596244 358912 596272
rect 303580 596232 303586 596244
rect 358906 596232 358912 596244
rect 358964 596232 358970 596284
rect 430666 596232 430672 596284
rect 430724 596272 430730 596284
rect 448514 596272 448520 596284
rect 430724 596244 448520 596272
rect 430724 596232 430730 596244
rect 448514 596232 448520 596244
rect 448572 596232 448578 596284
rect 39114 596164 39120 596216
rect 39172 596204 39178 596216
rect 55398 596204 55404 596216
rect 39172 596176 55404 596204
rect 39172 596164 39178 596176
rect 55398 596164 55404 596176
rect 55456 596164 55462 596216
rect 91002 596164 91008 596216
rect 91060 596204 91066 596216
rect 200758 596204 200764 596216
rect 91060 596176 200764 596204
rect 91060 596164 91066 596176
rect 200758 596164 200764 596176
rect 200816 596164 200822 596216
rect 255406 596164 255412 596216
rect 255464 596204 255470 596216
rect 273254 596204 273260 596216
rect 255464 596176 273260 596204
rect 255464 596164 255470 596176
rect 273254 596164 273260 596176
rect 273312 596164 273318 596216
rect 296346 596164 296352 596216
rect 296404 596204 296410 596216
rect 357802 596204 357808 596216
rect 296404 596176 357808 596204
rect 296404 596164 296410 596176
rect 357802 596164 357808 596176
rect 357860 596164 357866 596216
rect 399846 596164 399852 596216
rect 399904 596204 399910 596216
rect 415394 596204 415400 596216
rect 399904 596176 415400 596204
rect 399904 596164 399910 596176
rect 415394 596164 415400 596176
rect 415452 596164 415458 596216
rect 437474 596164 437480 596216
rect 437532 596204 437538 596216
rect 456794 596204 456800 596216
rect 437532 596176 456800 596204
rect 437532 596164 437538 596176
rect 456794 596164 456800 596176
rect 456852 596164 456858 596216
rect 216306 594736 216312 594788
rect 216364 594776 216370 594788
rect 249886 594776 249892 594788
rect 216364 594748 249892 594776
rect 216364 594736 216370 594748
rect 249886 594736 249892 594748
rect 249944 594736 249950 594788
rect 390186 594736 390192 594788
rect 390244 594776 390250 594788
rect 477494 594776 477500 594788
rect 390244 594748 477500 594776
rect 390244 594736 390250 594748
rect 477494 594736 477500 594748
rect 477552 594736 477558 594788
rect 218698 594668 218704 594720
rect 218756 594708 218762 594720
rect 253474 594708 253480 594720
rect 218756 594680 253480 594708
rect 218756 594668 218762 594680
rect 253474 594668 253480 594680
rect 253532 594668 253538 594720
rect 389910 594668 389916 594720
rect 389968 594708 389974 594720
rect 480254 594708 480260 594720
rect 389968 594680 480260 594708
rect 389968 594668 389974 594680
rect 480254 594668 480260 594680
rect 480312 594668 480318 594720
rect 217318 594600 217324 594652
rect 217376 594640 217382 594652
rect 252094 594640 252100 594652
rect 217376 594612 252100 594640
rect 217376 594600 217382 594612
rect 252094 594600 252100 594612
rect 252152 594600 252158 594652
rect 387518 594600 387524 594652
rect 387576 594640 387582 594652
rect 483014 594640 483020 594652
rect 387576 594612 483020 594640
rect 387576 594600 387582 594612
rect 483014 594600 483020 594612
rect 483072 594600 483078 594652
rect 214558 594532 214564 594584
rect 214616 594572 214622 594584
rect 255406 594572 255412 594584
rect 214616 594544 255412 594572
rect 214616 594532 214622 594544
rect 255406 594532 255412 594544
rect 255464 594532 255470 594584
rect 387150 594532 387156 594584
rect 387208 594572 387214 594584
rect 485774 594572 485780 594584
rect 387208 594544 485780 594572
rect 387208 594532 387214 594544
rect 485774 594532 485780 594544
rect 485832 594532 485838 594584
rect 214650 594464 214656 594516
rect 214708 594504 214714 594516
rect 259454 594504 259460 594516
rect 214708 594476 259460 594504
rect 214708 594464 214714 594476
rect 259454 594464 259460 594476
rect 259512 594464 259518 594516
rect 387334 594464 387340 594516
rect 387392 594504 387398 594516
rect 488534 594504 488540 594516
rect 387392 594476 488540 594504
rect 387392 594464 387398 594476
rect 488534 594464 488540 594476
rect 488592 594464 488598 594516
rect 214466 594396 214472 594448
rect 214524 594436 214530 594448
rect 259546 594436 259552 594448
rect 214524 594408 259552 594436
rect 214524 594396 214530 594408
rect 259546 594396 259552 594408
rect 259604 594396 259610 594448
rect 387610 594396 387616 594448
rect 387668 594436 387674 594448
rect 489914 594436 489920 594448
rect 387668 594408 489920 594436
rect 387668 594396 387674 594408
rect 489914 594396 489920 594408
rect 489972 594396 489978 594448
rect 219894 594328 219900 594380
rect 219952 594368 219958 594380
rect 285674 594368 285680 594380
rect 219952 594340 285680 594368
rect 219952 594328 219958 594340
rect 285674 594328 285680 594340
rect 285732 594328 285738 594380
rect 387426 594328 387432 594380
rect 387484 594368 387490 594380
rect 492674 594368 492680 594380
rect 387484 594340 492680 594368
rect 387484 594328 387490 594340
rect 492674 594328 492680 594340
rect 492732 594328 492738 594380
rect 212350 594260 212356 594312
rect 212408 594300 212414 594312
rect 280154 594300 280160 594312
rect 212408 594272 280160 594300
rect 212408 594260 212414 594272
rect 280154 594260 280160 594272
rect 280212 594260 280218 594312
rect 387242 594260 387248 594312
rect 387300 594300 387306 594312
rect 495434 594300 495440 594312
rect 387300 594272 495440 594300
rect 387300 594260 387306 594272
rect 495434 594260 495440 594272
rect 495492 594260 495498 594312
rect 36630 594192 36636 594244
rect 36688 594232 36694 594244
rect 71774 594232 71780 594244
rect 36688 594204 71780 594232
rect 36688 594192 36694 594204
rect 71774 594192 71780 594204
rect 71832 594192 71838 594244
rect 210970 594192 210976 594244
rect 211028 594232 211034 594244
rect 287054 594232 287060 594244
rect 211028 594204 287060 594232
rect 211028 594192 211034 594204
rect 287054 594192 287060 594204
rect 287112 594192 287118 594244
rect 387058 594192 387064 594244
rect 387116 594232 387122 594244
rect 498194 594232 498200 594244
rect 387116 594204 498200 594232
rect 387116 594192 387122 594204
rect 498194 594192 498200 594204
rect 498252 594192 498258 594244
rect 35802 594124 35808 594176
rect 35860 594164 35866 594176
rect 73154 594164 73160 594176
rect 35860 594136 73160 594164
rect 35860 594124 35866 594136
rect 73154 594124 73160 594136
rect 73212 594124 73218 594176
rect 215202 594124 215208 594176
rect 215260 594164 215266 594176
rect 292574 594164 292580 594176
rect 215260 594136 292580 594164
rect 215260 594124 215266 594136
rect 292574 594124 292580 594136
rect 292632 594124 292638 594176
rect 387702 594124 387708 594176
rect 387760 594164 387766 594176
rect 500954 594164 500960 594176
rect 387760 594136 500960 594164
rect 387760 594124 387766 594136
rect 500954 594124 500960 594136
rect 501012 594124 501018 594176
rect 36722 594056 36728 594108
rect 36780 594096 36786 594108
rect 76006 594096 76012 594108
rect 36780 594068 76012 594096
rect 36780 594056 36786 594068
rect 76006 594056 76012 594068
rect 76064 594056 76070 594108
rect 212442 594056 212448 594108
rect 212500 594096 212506 594108
rect 289814 594096 289820 594108
rect 212500 594068 289820 594096
rect 212500 594056 212506 594068
rect 289814 594056 289820 594068
rect 289872 594056 289878 594108
rect 386966 594056 386972 594108
rect 387024 594096 387030 594108
rect 502334 594096 502340 594108
rect 387024 594068 502340 594096
rect 387024 594056 387030 594068
rect 502334 594056 502340 594068
rect 502392 594056 502398 594108
rect 214374 593988 214380 594040
rect 214432 594028 214438 594040
rect 247126 594028 247132 594040
rect 214432 594000 247132 594028
rect 214432 593988 214438 594000
rect 247126 593988 247132 594000
rect 247184 593988 247190 594040
rect 390370 593988 390376 594040
rect 390428 594028 390434 594040
rect 474734 594028 474740 594040
rect 390428 594000 474740 594028
rect 390428 593988 390434 594000
rect 474734 593988 474740 594000
rect 474792 593988 474798 594040
rect 216490 593920 216496 593972
rect 216548 593960 216554 593972
rect 248414 593960 248420 593972
rect 216548 593932 248420 593960
rect 216548 593920 216554 593932
rect 248414 593920 248420 593932
rect 248472 593920 248478 593972
rect 390002 593920 390008 593972
rect 390060 593960 390066 593972
rect 473354 593960 473360 593972
rect 390060 593932 473360 593960
rect 390060 593920 390066 593932
rect 473354 593920 473360 593932
rect 473412 593920 473418 593972
rect 219342 593852 219348 593904
rect 219400 593892 219406 593904
rect 252186 593892 252192 593904
rect 219400 593864 252192 593892
rect 219400 593852 219406 593864
rect 252186 593852 252192 593864
rect 252244 593852 252250 593904
rect 395062 593852 395068 593904
rect 395120 593892 395126 593904
rect 438854 593892 438860 593904
rect 395120 593864 438860 593892
rect 395120 593852 395126 593864
rect 438854 593852 438860 593864
rect 438912 593852 438918 593904
rect 398006 591948 398012 592000
rect 398064 591988 398070 592000
rect 426434 591988 426440 592000
rect 398064 591960 426440 591988
rect 398064 591948 398070 591960
rect 426434 591948 426440 591960
rect 426492 591948 426498 592000
rect 399294 591880 399300 591932
rect 399352 591920 399358 591932
rect 429194 591920 429200 591932
rect 399352 591892 429200 591920
rect 399352 591880 399358 591892
rect 429194 591880 429200 591892
rect 429252 591880 429258 591932
rect 397914 591812 397920 591864
rect 397972 591852 397978 591864
rect 427998 591852 428004 591864
rect 397972 591824 428004 591852
rect 397972 591812 397978 591824
rect 427998 591812 428004 591824
rect 428056 591812 428062 591864
rect 398190 591744 398196 591796
rect 398248 591784 398254 591796
rect 430666 591784 430672 591796
rect 398248 591756 430672 591784
rect 398248 591744 398254 591756
rect 430666 591744 430672 591756
rect 430724 591744 430730 591796
rect 399202 591676 399208 591728
rect 399260 591716 399266 591728
rect 431954 591716 431960 591728
rect 399260 591688 431960 591716
rect 399260 591676 399266 591688
rect 431954 591676 431960 591688
rect 432012 591676 432018 591728
rect 399386 591608 399392 591660
rect 399444 591648 399450 591660
rect 433426 591648 433432 591660
rect 399444 591620 433432 591648
rect 399444 591608 399450 591620
rect 433426 591608 433432 591620
rect 433484 591608 433490 591660
rect 395798 591540 395804 591592
rect 395856 591580 395862 591592
rect 437474 591580 437480 591592
rect 395856 591552 437480 591580
rect 395856 591540 395862 591552
rect 437474 591540 437480 591552
rect 437532 591540 437538 591592
rect 395154 591472 395160 591524
rect 395212 591512 395218 591524
rect 440326 591512 440332 591524
rect 395212 591484 440332 591512
rect 395212 591472 395218 591484
rect 440326 591472 440332 591484
rect 440384 591472 440390 591524
rect 384390 591404 384396 591456
rect 384448 591444 384454 591456
rect 445754 591444 445760 591456
rect 384448 591416 445760 591444
rect 384448 591404 384454 591416
rect 445754 591404 445760 591416
rect 445812 591404 445818 591456
rect 384298 591336 384304 591388
rect 384356 591376 384362 591388
rect 447134 591376 447140 591388
rect 384356 591348 447140 591376
rect 384356 591336 384362 591348
rect 447134 591336 447140 591348
rect 447192 591336 447198 591388
rect 384482 591268 384488 591320
rect 384540 591308 384546 591320
rect 449894 591308 449900 591320
rect 384540 591280 449900 591308
rect 384540 591268 384546 591280
rect 449894 591268 449900 591280
rect 449952 591268 449958 591320
rect 188338 590656 188344 590708
rect 188396 590696 188402 590708
rect 579614 590696 579620 590708
rect 188396 590668 579620 590696
rect 188396 590656 188402 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 38470 585760 38476 585812
rect 38528 585800 38534 585812
rect 217134 585800 217140 585812
rect 38528 585772 217140 585800
rect 38528 585760 38534 585772
rect 217134 585760 217140 585772
rect 217192 585760 217198 585812
rect 37734 585148 37740 585200
rect 37792 585188 37798 585200
rect 38470 585188 38476 585200
rect 37792 585160 38476 585188
rect 37792 585148 37798 585160
rect 38470 585148 38476 585160
rect 38528 585148 38534 585200
rect 2774 579912 2780 579964
rect 2832 579952 2838 579964
rect 4890 579952 4896 579964
rect 2832 579924 4896 579952
rect 2832 579912 2838 579924
rect 4890 579912 4896 579924
rect 4948 579912 4954 579964
rect 193858 576852 193864 576904
rect 193916 576892 193922 576904
rect 579614 576892 579620 576904
rect 193916 576864 579620 576892
rect 193916 576852 193922 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 170858 567128 170864 567180
rect 170916 567168 170922 567180
rect 213914 567168 213920 567180
rect 170916 567140 213920 567168
rect 170916 567128 170922 567140
rect 213914 567128 213920 567140
rect 213972 567128 213978 567180
rect 351086 567128 351092 567180
rect 351144 567168 351150 567180
rect 394694 567168 394700 567180
rect 351144 567140 394700 567168
rect 351144 567128 351150 567140
rect 394694 567128 394700 567140
rect 394752 567128 394758 567180
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 35158 565876 35164 565888
rect 3476 565848 35164 565876
rect 3476 565836 3482 565848
rect 35158 565836 35164 565848
rect 35216 565836 35222 565888
rect 530946 565836 530952 565888
rect 531004 565876 531010 565888
rect 536834 565876 536840 565888
rect 531004 565848 536840 565876
rect 531004 565836 531010 565848
rect 536834 565836 536840 565848
rect 536892 565836 536898 565888
rect 142062 565700 142068 565752
rect 142120 565740 142126 565752
rect 204070 565740 204076 565752
rect 142120 565712 204076 565740
rect 142120 565700 142126 565712
rect 204070 565700 204076 565712
rect 204128 565700 204134 565752
rect 136542 565632 136548 565684
rect 136600 565672 136606 565684
rect 203886 565672 203892 565684
rect 136600 565644 203892 565672
rect 136600 565632 136606 565644
rect 203886 565632 203892 565644
rect 203944 565632 203950 565684
rect 133782 565564 133788 565616
rect 133840 565604 133846 565616
rect 203794 565604 203800 565616
rect 133840 565576 203800 565604
rect 133840 565564 133846 565576
rect 203794 565564 203800 565576
rect 203852 565564 203858 565616
rect 131022 565496 131028 565548
rect 131080 565536 131086 565548
rect 203702 565536 203708 565548
rect 131080 565508 203708 565536
rect 131080 565496 131086 565508
rect 203702 565496 203708 565508
rect 203760 565496 203766 565548
rect 88242 565428 88248 565480
rect 88300 565468 88306 565480
rect 200942 565468 200948 565480
rect 88300 565440 200948 565468
rect 88300 565428 88306 565440
rect 200942 565428 200948 565440
rect 201000 565428 201006 565480
rect 86862 565360 86868 565412
rect 86920 565400 86926 565412
rect 200850 565400 200856 565412
rect 86920 565372 200856 565400
rect 86920 565360 86926 565372
rect 200850 565360 200856 565372
rect 200908 565360 200914 565412
rect 84102 565292 84108 565344
rect 84160 565332 84166 565344
rect 201034 565332 201040 565344
rect 84160 565304 201040 565332
rect 84160 565292 84166 565304
rect 201034 565292 201040 565304
rect 201092 565292 201098 565344
rect 81342 565224 81348 565276
rect 81400 565264 81406 565276
rect 203978 565264 203984 565276
rect 81400 565236 203984 565264
rect 81400 565224 81406 565236
rect 203978 565224 203984 565236
rect 204036 565224 204042 565276
rect 78582 565156 78588 565208
rect 78640 565196 78646 565208
rect 203610 565196 203616 565208
rect 78640 565168 203616 565196
rect 78640 565156 78646 565168
rect 203610 565156 203616 565168
rect 203668 565156 203674 565208
rect 77202 565088 77208 565140
rect 77260 565128 77266 565140
rect 203518 565128 203524 565140
rect 77260 565100 203524 565128
rect 77260 565088 77266 565100
rect 203518 565088 203524 565100
rect 203576 565088 203582 565140
rect 214926 563728 214932 563780
rect 214984 563768 214990 563780
rect 249794 563768 249800 563780
rect 214984 563740 249800 563768
rect 214984 563728 214990 563740
rect 249794 563728 249800 563740
rect 249852 563728 249858 563780
rect 37826 563660 37832 563712
rect 37884 563700 37890 563712
rect 217226 563700 217232 563712
rect 37884 563672 217232 563700
rect 37884 563660 37890 563672
rect 217226 563660 217232 563672
rect 217284 563660 217290 563712
rect 39022 563252 39028 563304
rect 39080 563292 39086 563304
rect 40034 563292 40040 563304
rect 39080 563264 40040 563292
rect 39080 563252 39086 563264
rect 40034 563252 40040 563264
rect 40092 563252 40098 563304
rect 537662 563048 537668 563100
rect 537720 563088 537726 563100
rect 579890 563088 579896 563100
rect 537720 563060 579896 563088
rect 537720 563048 537726 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 25590 553432 25596 553444
rect 3476 553404 25596 553432
rect 3476 553392 3482 553404
rect 25590 553392 25596 553404
rect 25648 553392 25654 553444
rect 544378 536800 544384 536852
rect 544436 536840 544442 536852
rect 580166 536840 580172 536852
rect 544436 536812 580172 536840
rect 544436 536800 544442 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527824 3424 527876
rect 3476 527864 3482 527876
rect 8938 527864 8944 527876
rect 3476 527836 8944 527864
rect 3476 527824 3482 527836
rect 8938 527824 8944 527836
rect 8996 527824 9002 527876
rect 541618 524424 541624 524476
rect 541676 524464 541682 524476
rect 580166 524464 580172 524476
rect 541676 524436 580172 524464
rect 541676 524424 541682 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 537570 510620 537576 510672
rect 537628 510660 537634 510672
rect 580166 510660 580172 510672
rect 537628 510632 580172 510660
rect 537628 510620 537634 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 14458 501004 14464 501016
rect 3108 500976 14464 501004
rect 3108 500964 3114 500976
rect 14458 500964 14464 500976
rect 14516 500964 14522 501016
rect 374638 487772 374644 487824
rect 374696 487812 374702 487824
rect 397178 487812 397184 487824
rect 374696 487784 397184 487812
rect 374696 487772 374702 487784
rect 397178 487772 397184 487784
rect 397236 487772 397242 487824
rect 39022 485256 39028 485308
rect 39080 485296 39086 485308
rect 39666 485296 39672 485308
rect 39080 485268 39672 485296
rect 39080 485256 39086 485268
rect 39666 485256 39672 485268
rect 39724 485256 39730 485308
rect 39758 485256 39764 485308
rect 39816 485256 39822 485308
rect 39776 485104 39804 485256
rect 39758 485052 39764 485104
rect 39816 485052 39822 485104
rect 38930 484916 38936 484968
rect 38988 484956 38994 484968
rect 39942 484956 39948 484968
rect 38988 484928 39948 484956
rect 38988 484916 38994 484928
rect 39942 484916 39948 484928
rect 40000 484916 40006 484968
rect 540238 484372 540244 484424
rect 540296 484412 540302 484424
rect 580166 484412 580172 484424
rect 540296 484384 580172 484412
rect 540296 484372 540302 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 38102 480020 38108 480072
rect 38160 480060 38166 480072
rect 217594 480060 217600 480072
rect 38160 480032 217600 480060
rect 38160 480020 38166 480032
rect 217594 480020 217600 480032
rect 217652 480020 217658 480072
rect 38286 479952 38292 480004
rect 38344 479992 38350 480004
rect 216858 479992 216864 480004
rect 38344 479964 216864 479992
rect 38344 479952 38350 479964
rect 216858 479952 216864 479964
rect 216916 479952 216922 480004
rect 38562 479884 38568 479936
rect 38620 479924 38626 479936
rect 216674 479924 216680 479936
rect 38620 479896 216680 479924
rect 38620 479884 38626 479896
rect 216674 479884 216680 479896
rect 216732 479884 216738 479936
rect 38010 479816 38016 479868
rect 38068 479856 38074 479868
rect 217134 479856 217140 479868
rect 38068 479828 217140 479856
rect 38068 479816 38074 479828
rect 217134 479816 217140 479828
rect 217192 479816 217198 479868
rect 37826 479748 37832 479800
rect 37884 479788 37890 479800
rect 217410 479788 217416 479800
rect 37884 479760 217416 479788
rect 37884 479748 37890 479760
rect 217410 479748 217416 479760
rect 217468 479748 217474 479800
rect 216858 479476 216864 479528
rect 216916 479516 216922 479528
rect 217502 479516 217508 479528
rect 216916 479488 217508 479516
rect 216916 479476 216922 479488
rect 217502 479476 217508 479488
rect 217560 479476 217566 479528
rect 216674 479340 216680 479392
rect 216732 479380 216738 479392
rect 217778 479380 217784 479392
rect 216732 479352 217784 479380
rect 216732 479340 216738 479352
rect 217778 479340 217784 479352
rect 217836 479340 217842 479392
rect 218330 478972 218336 478984
rect 200086 478944 218336 478972
rect 39114 478864 39120 478916
rect 39172 478904 39178 478916
rect 56042 478904 56048 478916
rect 39172 478876 56048 478904
rect 39172 478864 39178 478876
rect 56042 478864 56048 478876
rect 56100 478904 56106 478916
rect 200086 478904 200114 478944
rect 218330 478932 218336 478944
rect 218388 478972 218394 478984
rect 218388 478944 219434 478972
rect 218388 478932 218394 478944
rect 56100 478876 200114 478904
rect 56100 478864 56106 478876
rect 217226 478864 217232 478916
rect 217284 478904 217290 478916
rect 217594 478904 217600 478916
rect 217284 478876 217600 478904
rect 217284 478864 217290 478876
rect 217594 478864 217600 478876
rect 217652 478864 217658 478916
rect 219406 478904 219434 478944
rect 219710 478904 219716 478916
rect 219406 478876 219716 478904
rect 219710 478864 219716 478876
rect 219768 478904 219774 478916
rect 235994 478904 236000 478916
rect 219768 478876 236000 478904
rect 219768 478864 219774 478876
rect 235994 478864 236000 478876
rect 236052 478864 236058 478916
rect 36630 478592 36636 478644
rect 36688 478632 36694 478644
rect 72326 478632 72332 478644
rect 36688 478604 72332 478632
rect 36688 478592 36694 478604
rect 72326 478592 72332 478604
rect 72384 478632 72390 478644
rect 73798 478632 73804 478644
rect 72384 478604 73804 478632
rect 72384 478592 72390 478604
rect 73798 478592 73804 478604
rect 73856 478592 73862 478644
rect 39206 478524 39212 478576
rect 39264 478564 39270 478576
rect 74626 478564 74632 478576
rect 39264 478536 74632 478564
rect 39264 478524 39270 478536
rect 74626 478524 74632 478536
rect 74684 478564 74690 478576
rect 77202 478564 77208 478576
rect 74684 478536 77208 478564
rect 74684 478524 74690 478536
rect 77202 478524 77208 478536
rect 77260 478524 77266 478576
rect 398374 478524 398380 478576
rect 398432 478564 398438 478576
rect 425514 478564 425520 478576
rect 398432 478536 425520 478564
rect 398432 478524 398438 478536
rect 425514 478524 425520 478536
rect 425572 478524 425578 478576
rect 35802 478456 35808 478508
rect 35860 478496 35866 478508
rect 73154 478496 73160 478508
rect 35860 478468 73160 478496
rect 35860 478456 35866 478468
rect 73154 478456 73160 478468
rect 73212 478456 73218 478508
rect 399570 478456 399576 478508
rect 399628 478496 399634 478508
rect 426618 478496 426624 478508
rect 399628 478468 426624 478496
rect 399628 478456 399634 478468
rect 426618 478456 426624 478468
rect 426676 478456 426682 478508
rect 37918 478388 37924 478440
rect 37976 478428 37982 478440
rect 76926 478428 76932 478440
rect 37976 478400 76932 478428
rect 37976 478388 37982 478400
rect 76926 478388 76932 478400
rect 76984 478428 76990 478440
rect 78582 478428 78588 478440
rect 76984 478400 78588 478428
rect 76984 478388 76990 478400
rect 78582 478388 78588 478400
rect 78640 478388 78646 478440
rect 398006 478388 398012 478440
rect 398064 478428 398070 478440
rect 427814 478428 427820 478440
rect 398064 478400 427820 478428
rect 398064 478388 398070 478400
rect 427814 478388 427820 478400
rect 427872 478388 427878 478440
rect 36722 478320 36728 478372
rect 36780 478360 36786 478372
rect 75822 478360 75828 478372
rect 36780 478332 75828 478360
rect 36780 478320 36786 478332
rect 75822 478320 75828 478332
rect 75880 478360 75886 478372
rect 78214 478360 78220 478372
rect 75880 478332 78220 478360
rect 75880 478320 75886 478332
rect 78214 478320 78220 478332
rect 78272 478320 78278 478372
rect 399294 478320 399300 478372
rect 399352 478360 399358 478372
rect 430114 478360 430120 478372
rect 399352 478332 430120 478360
rect 399352 478320 399358 478332
rect 430114 478320 430120 478332
rect 430172 478360 430178 478372
rect 430574 478360 430580 478372
rect 430172 478332 430580 478360
rect 430172 478320 430178 478332
rect 430574 478320 430580 478332
rect 430632 478320 430638 478372
rect 36906 478252 36912 478304
rect 36964 478292 36970 478304
rect 78122 478292 78128 478304
rect 36964 478264 78128 478292
rect 36964 478252 36970 478264
rect 78122 478252 78128 478264
rect 78180 478252 78186 478304
rect 397914 478252 397920 478304
rect 397972 478292 397978 478304
rect 428550 478292 428556 478304
rect 397972 478264 428556 478292
rect 397972 478252 397978 478264
rect 428550 478252 428556 478264
rect 428608 478292 428614 478304
rect 430022 478292 430028 478304
rect 428608 478264 430028 478292
rect 428608 478252 428614 478264
rect 430022 478252 430028 478264
rect 430080 478252 430086 478304
rect 36998 478184 37004 478236
rect 37056 478224 37062 478236
rect 79502 478224 79508 478236
rect 37056 478196 79508 478224
rect 37056 478184 37062 478196
rect 79502 478184 79508 478196
rect 79560 478184 79566 478236
rect 398190 478184 398196 478236
rect 398248 478224 398254 478236
rect 431310 478224 431316 478236
rect 398248 478196 431316 478224
rect 398248 478184 398254 478196
rect 431310 478184 431316 478196
rect 431368 478224 431374 478236
rect 433242 478224 433248 478236
rect 431368 478196 433248 478224
rect 431368 478184 431374 478196
rect 433242 478184 433248 478196
rect 433300 478184 433306 478236
rect 36814 478116 36820 478168
rect 36872 478156 36878 478168
rect 80606 478156 80612 478168
rect 36872 478128 80612 478156
rect 36872 478116 36878 478128
rect 80606 478116 80612 478128
rect 80664 478156 80670 478168
rect 82722 478156 82728 478168
rect 80664 478128 82728 478156
rect 80664 478116 80670 478128
rect 82722 478116 82728 478128
rect 82780 478116 82786 478168
rect 399202 478116 399208 478168
rect 399260 478156 399266 478168
rect 432506 478156 432512 478168
rect 399260 478128 432512 478156
rect 399260 478116 399266 478128
rect 432506 478116 432512 478128
rect 432564 478156 432570 478168
rect 434622 478156 434628 478168
rect 432564 478128 434628 478156
rect 432564 478116 432570 478128
rect 434622 478116 434628 478128
rect 434680 478116 434686 478168
rect 394326 477912 394332 477964
rect 394384 477952 394390 477964
rect 398374 477952 398380 477964
rect 394384 477924 398380 477952
rect 394384 477912 394390 477924
rect 398374 477912 398380 477924
rect 398432 477912 398438 477964
rect 394418 477844 394424 477896
rect 394476 477884 394482 477896
rect 399570 477884 399576 477896
rect 394476 477856 399576 477884
rect 394476 477844 394482 477856
rect 399570 477844 399576 477856
rect 399628 477844 399634 477896
rect 397270 477776 397276 477828
rect 397328 477816 397334 477828
rect 399294 477816 399300 477828
rect 397328 477788 399300 477816
rect 397328 477776 397334 477788
rect 399294 477776 399300 477788
rect 399352 477776 399358 477828
rect 394510 477708 394516 477760
rect 394568 477748 394574 477760
rect 398006 477748 398012 477760
rect 394568 477720 398012 477748
rect 394568 477708 394574 477720
rect 398006 477708 398012 477720
rect 398064 477708 398070 477760
rect 398282 477708 398288 477760
rect 398340 477748 398346 477760
rect 400122 477748 400128 477760
rect 398340 477720 400128 477748
rect 398340 477708 398346 477720
rect 400122 477708 400128 477720
rect 400180 477708 400186 477760
rect 394602 477640 394608 477692
rect 394660 477680 394666 477692
rect 397914 477680 397920 477692
rect 394660 477652 397920 477680
rect 394660 477640 394666 477652
rect 397914 477640 397920 477652
rect 397972 477640 397978 477692
rect 398466 477640 398472 477692
rect 398524 477680 398530 477692
rect 424134 477680 424140 477692
rect 398524 477652 424140 477680
rect 398524 477640 398530 477652
rect 424134 477640 424140 477652
rect 424192 477680 424198 477692
rect 426158 477680 426164 477692
rect 424192 477652 426164 477680
rect 424192 477640 424198 477652
rect 426158 477640 426164 477652
rect 426216 477640 426222 477692
rect 397178 477572 397184 477624
rect 397236 477612 397242 477624
rect 398098 477612 398104 477624
rect 397236 477584 398104 477612
rect 397236 477572 397242 477584
rect 398098 477572 398104 477584
rect 398156 477572 398162 477624
rect 399018 477572 399024 477624
rect 399076 477612 399082 477624
rect 399478 477612 399484 477624
rect 399076 477584 399484 477612
rect 399076 477572 399082 477584
rect 399478 477572 399484 477584
rect 399536 477612 399542 477624
rect 436002 477612 436008 477624
rect 399536 477584 436008 477612
rect 399536 477572 399542 477584
rect 397362 477504 397368 477556
rect 397420 477544 397426 477556
rect 398190 477544 398196 477556
rect 397420 477516 398196 477544
rect 397420 477504 397426 477516
rect 398190 477504 398196 477516
rect 398248 477504 398254 477556
rect 398742 477504 398748 477556
rect 398800 477544 398806 477556
rect 399202 477544 399208 477556
rect 398800 477516 399208 477544
rect 398800 477504 398806 477516
rect 399202 477504 399208 477516
rect 399260 477504 399266 477556
rect 399386 477504 399392 477556
rect 399444 477544 399450 477556
rect 434438 477544 434444 477556
rect 399444 477516 434444 477544
rect 399444 477504 399450 477516
rect 433444 477488 433472 477516
rect 434438 477504 434444 477516
rect 434496 477504 434502 477556
rect 434548 477488 434576 477584
rect 436002 477572 436008 477584
rect 436060 477572 436066 477624
rect 37090 477436 37096 477488
rect 37148 477476 37154 477488
rect 70854 477476 70860 477488
rect 37148 477448 70860 477476
rect 37148 477436 37154 477448
rect 70854 477436 70860 477448
rect 70912 477436 70918 477488
rect 86954 477436 86960 477488
rect 87012 477476 87018 477488
rect 87598 477476 87604 477488
rect 87012 477448 87604 477476
rect 87012 477436 87018 477448
rect 87598 477436 87604 477448
rect 87656 477476 87662 477488
rect 216490 477476 216496 477488
rect 87656 477448 216496 477476
rect 87656 477436 87662 477448
rect 216490 477436 216496 477448
rect 216548 477436 216554 477488
rect 217042 477436 217048 477488
rect 217100 477476 217106 477488
rect 217318 477476 217324 477488
rect 217100 477448 217324 477476
rect 217100 477436 217106 477448
rect 217318 477436 217324 477448
rect 217376 477476 217382 477488
rect 252370 477476 252376 477488
rect 217376 477448 252376 477476
rect 217376 477436 217382 477448
rect 252370 477436 252376 477448
rect 252428 477436 252434 477488
rect 252462 477436 252468 477488
rect 252520 477476 252526 477488
rect 269114 477476 269120 477488
rect 252520 477448 269120 477476
rect 252520 477436 252526 477448
rect 269114 477436 269120 477448
rect 269172 477436 269178 477488
rect 433426 477436 433432 477488
rect 433484 477436 433490 477488
rect 434530 477436 434536 477488
rect 434588 477436 434594 477488
rect 37182 477368 37188 477420
rect 37240 477408 37246 477420
rect 70210 477408 70216 477420
rect 37240 477380 70216 477408
rect 37240 477368 37246 477380
rect 70210 477368 70216 477380
rect 70268 477368 70274 477420
rect 85574 477368 85580 477420
rect 85632 477408 85638 477420
rect 86310 477408 86316 477420
rect 85632 477380 86316 477408
rect 85632 477368 85638 477380
rect 86310 477368 86316 477380
rect 86368 477408 86374 477420
rect 214374 477408 214380 477420
rect 86368 477380 214380 477408
rect 86368 477368 86374 477380
rect 214374 477368 214380 477380
rect 214432 477368 214438 477420
rect 214558 477368 214564 477420
rect 214616 477408 214622 477420
rect 255314 477408 255320 477420
rect 214616 477380 255320 477408
rect 214616 477368 214622 477380
rect 255314 477368 255320 477380
rect 255372 477368 255378 477420
rect 260834 477368 260840 477420
rect 260892 477408 260898 477420
rect 278774 477408 278780 477420
rect 260892 477380 278780 477408
rect 260892 477368 260898 477380
rect 278774 477368 278780 477380
rect 278832 477368 278838 477420
rect 433242 477368 433248 477420
rect 433300 477408 433306 477420
rect 448514 477408 448520 477420
rect 433300 477380 448520 477408
rect 433300 477368 433306 477380
rect 448514 477368 448520 477380
rect 448572 477368 448578 477420
rect 37642 477300 37648 477352
rect 37700 477340 37706 477352
rect 67634 477340 67640 477352
rect 37700 477312 67640 477340
rect 37700 477300 37706 477312
rect 67634 477300 67640 477312
rect 67692 477340 67698 477352
rect 67692 477312 74534 477340
rect 67692 477300 67698 477312
rect 39298 477232 39304 477284
rect 39356 477272 39362 477284
rect 68738 477272 68744 477284
rect 39356 477244 68744 477272
rect 39356 477232 39362 477244
rect 68738 477232 68744 477244
rect 68796 477272 68802 477284
rect 68796 477244 69428 477272
rect 68796 477232 68802 477244
rect 39390 477164 39396 477216
rect 39448 477204 39454 477216
rect 66530 477204 66536 477216
rect 39448 477176 66536 477204
rect 39448 477164 39454 477176
rect 66530 477164 66536 477176
rect 66588 477204 66594 477216
rect 67542 477204 67548 477216
rect 66588 477176 67548 477204
rect 66588 477164 66594 477176
rect 67542 477164 67548 477176
rect 67600 477164 67606 477216
rect 38378 477096 38384 477148
rect 38436 477136 38442 477148
rect 64874 477136 64880 477148
rect 38436 477108 64880 477136
rect 38436 477096 38442 477108
rect 64874 477096 64880 477108
rect 64932 477096 64938 477148
rect 69400 477136 69428 477244
rect 74506 477204 74534 477312
rect 78582 477300 78588 477352
rect 78640 477340 78646 477352
rect 95786 477340 95792 477352
rect 78640 477312 95792 477340
rect 78640 477300 78646 477312
rect 95786 477300 95792 477312
rect 95844 477340 95850 477352
rect 96522 477340 96528 477352
rect 95844 477312 96528 477340
rect 95844 477300 95850 477312
rect 96522 477300 96528 477312
rect 96580 477300 96586 477352
rect 214742 477340 214748 477352
rect 103486 477312 214748 477340
rect 78122 477232 78128 477284
rect 78180 477272 78186 477284
rect 96982 477272 96988 477284
rect 78180 477244 96988 477272
rect 78180 477232 78186 477244
rect 96982 477232 96988 477244
rect 97040 477272 97046 477284
rect 103486 477272 103514 477312
rect 214742 477300 214748 477312
rect 214800 477300 214806 477352
rect 215110 477300 215116 477352
rect 215168 477340 215174 477352
rect 245930 477340 245936 477352
rect 215168 477312 245936 477340
rect 215168 477300 215174 477312
rect 245930 477300 245936 477312
rect 245988 477300 245994 477352
rect 247126 477300 247132 477352
rect 247184 477340 247190 477352
rect 266354 477340 266360 477352
rect 247184 477312 266360 477340
rect 247184 477300 247190 477312
rect 266354 477300 266360 477312
rect 266412 477300 266418 477352
rect 436002 477300 436008 477352
rect 436060 477340 436066 477352
rect 452654 477340 452660 477352
rect 436060 477312 452660 477340
rect 436060 477300 436066 477312
rect 452654 477300 452660 477312
rect 452712 477300 452718 477352
rect 97040 477244 103514 477272
rect 97040 477232 97046 477244
rect 214834 477232 214840 477284
rect 214892 477272 214898 477284
rect 245470 477272 245476 477284
rect 214892 477244 245476 477272
rect 214892 477232 214898 477244
rect 245470 477232 245476 477244
rect 245528 477272 245534 477284
rect 263594 477272 263600 477284
rect 245528 477244 263600 477272
rect 245528 477232 245534 477244
rect 263594 477232 263600 477244
rect 263652 477232 263658 477284
rect 263686 477232 263692 477284
rect 263744 477272 263750 477284
rect 277670 477272 277676 477284
rect 263744 477244 277676 477272
rect 263744 477232 263750 477244
rect 277670 477232 277676 477244
rect 277728 477232 277734 477284
rect 430022 477232 430028 477284
rect 430080 477272 430086 477284
rect 447134 477272 447140 477284
rect 430080 477244 447140 477272
rect 430080 477232 430086 477244
rect 447134 477232 447140 477244
rect 447192 477232 447198 477284
rect 85574 477204 85580 477216
rect 74506 477176 85580 477204
rect 85574 477164 85580 477176
rect 85632 477164 85638 477216
rect 207014 477164 207020 477216
rect 207072 477204 207078 477216
rect 208302 477204 208308 477216
rect 207072 477176 208308 477204
rect 207072 477164 207078 477176
rect 208302 477164 208308 477176
rect 208360 477204 208366 477216
rect 217042 477204 217048 477216
rect 208360 477176 217048 477204
rect 208360 477164 208366 477176
rect 217042 477164 217048 477176
rect 217100 477164 217106 477216
rect 219342 477164 219348 477216
rect 219400 477204 219406 477216
rect 251266 477204 251272 477216
rect 219400 477176 251272 477204
rect 219400 477164 219406 477176
rect 251266 477164 251272 477176
rect 251324 477204 251330 477216
rect 252462 477204 252468 477216
rect 251324 477176 252468 477204
rect 251324 477164 251330 477176
rect 252462 477164 252468 477176
rect 252520 477164 252526 477216
rect 259362 477164 259368 477216
rect 259420 477204 259426 477216
rect 276014 477204 276020 477216
rect 259420 477176 276020 477204
rect 259420 477164 259426 477176
rect 276014 477164 276020 477176
rect 276072 477164 276078 477216
rect 399662 477164 399668 477216
rect 399720 477204 399726 477216
rect 416774 477204 416780 477216
rect 399720 477176 416780 477204
rect 399720 477164 399726 477176
rect 416774 477164 416780 477176
rect 416832 477164 416838 477216
rect 430574 477164 430580 477216
rect 430632 477204 430638 477216
rect 448514 477204 448520 477216
rect 430632 477176 448520 477204
rect 430632 477164 430638 477176
rect 448514 477164 448520 477176
rect 448572 477164 448578 477216
rect 69400 477108 74534 477136
rect 39758 477028 39764 477080
rect 39816 477068 39822 477080
rect 63494 477068 63500 477080
rect 39816 477040 63500 477068
rect 39816 477028 39822 477040
rect 63494 477028 63500 477040
rect 63552 477028 63558 477080
rect 74506 477068 74534 477108
rect 77202 477096 77208 477148
rect 77260 477136 77266 477148
rect 93026 477136 93032 477148
rect 77260 477108 93032 477136
rect 77260 477096 77266 477108
rect 93026 477096 93032 477108
rect 93084 477096 93090 477148
rect 216398 477096 216404 477148
rect 216456 477136 216462 477148
rect 250070 477136 250076 477148
rect 216456 477108 250076 477136
rect 216456 477096 216462 477108
rect 250070 477096 250076 477108
rect 250128 477136 250134 477148
rect 251082 477136 251088 477148
rect 250128 477108 251088 477136
rect 250128 477096 250134 477108
rect 251082 477096 251088 477108
rect 251140 477096 251146 477148
rect 255314 477096 255320 477148
rect 255372 477136 255378 477148
rect 273254 477136 273260 477148
rect 255372 477108 273260 477136
rect 255372 477096 255378 477108
rect 273254 477096 273260 477108
rect 273312 477096 273318 477148
rect 399846 477096 399852 477148
rect 399904 477136 399910 477148
rect 415394 477136 415400 477148
rect 399904 477108 415400 477136
rect 399904 477096 399910 477108
rect 415394 477096 415400 477108
rect 415452 477096 415458 477148
rect 427722 477096 427728 477148
rect 427780 477136 427786 477148
rect 445754 477136 445760 477148
rect 427780 477108 445760 477136
rect 427780 477096 427786 477108
rect 445754 477096 445760 477108
rect 445812 477096 445818 477148
rect 86954 477068 86960 477080
rect 74506 477040 86960 477068
rect 86954 477028 86960 477040
rect 87012 477028 87018 477080
rect 96522 477028 96528 477080
rect 96580 477068 96586 477080
rect 215018 477068 215024 477080
rect 96580 477040 215024 477068
rect 96580 477028 96586 477040
rect 215018 477028 215024 477040
rect 215076 477068 215082 477080
rect 256970 477068 256976 477080
rect 215076 477040 256976 477068
rect 215076 477028 215082 477040
rect 256970 477028 256976 477040
rect 257028 477068 257034 477080
rect 274634 477068 274640 477080
rect 257028 477040 274640 477068
rect 257028 477028 257034 477040
rect 274634 477028 274640 477040
rect 274692 477028 274698 477080
rect 399938 477028 399944 477080
rect 399996 477068 400002 477080
rect 419534 477068 419540 477080
rect 399996 477040 419540 477068
rect 399996 477028 400002 477040
rect 419534 477028 419540 477040
rect 419592 477028 419598 477080
rect 426618 477028 426624 477080
rect 426676 477068 426682 477080
rect 444374 477068 444380 477080
rect 426676 477040 444380 477068
rect 426676 477028 426682 477040
rect 444374 477028 444380 477040
rect 444432 477028 444438 477080
rect 445662 477028 445668 477080
rect 445720 477068 445726 477080
rect 458174 477068 458180 477080
rect 445720 477040 458180 477068
rect 445720 477028 445726 477040
rect 458174 477028 458180 477040
rect 458232 477028 458238 477080
rect 39482 476960 39488 477012
rect 39540 477000 39546 477012
rect 63218 477000 63224 477012
rect 39540 476972 63224 477000
rect 39540 476960 39546 476972
rect 63218 476960 63224 476972
rect 63276 477000 63282 477012
rect 63276 476972 64874 477000
rect 63276 476960 63282 476972
rect 39574 476892 39580 476944
rect 39632 476932 39638 476944
rect 60734 476932 60740 476944
rect 39632 476904 60740 476932
rect 39632 476892 39638 476904
rect 60734 476892 60740 476904
rect 60792 476892 60798 476944
rect 39022 476824 39028 476876
rect 39080 476864 39086 476876
rect 59446 476864 59452 476876
rect 39080 476836 59452 476864
rect 39080 476824 39086 476836
rect 59446 476824 59452 476836
rect 59504 476824 59510 476876
rect 64846 476864 64874 476972
rect 70854 476960 70860 477012
rect 70912 477000 70918 477012
rect 89714 477000 89720 477012
rect 70912 476972 89720 477000
rect 70912 476960 70918 476972
rect 89714 476960 89720 476972
rect 89772 476960 89778 477012
rect 217962 476960 217968 477012
rect 218020 477000 218026 477012
rect 218790 477000 218796 477012
rect 218020 476972 218796 477000
rect 218020 476960 218026 476972
rect 218790 476960 218796 476972
rect 218848 477000 218854 477012
rect 244274 477000 244280 477012
rect 218848 476972 244280 477000
rect 218848 476960 218854 476972
rect 244274 476960 244280 476972
rect 244332 476960 244338 477012
rect 252370 476960 252376 477012
rect 252428 477000 252434 477012
rect 270494 477000 270500 477012
rect 252428 476972 270500 477000
rect 252428 476960 252434 476972
rect 270494 476960 270500 476972
rect 270552 476960 270558 477012
rect 399478 476960 399484 477012
rect 399536 477000 399542 477012
rect 400122 477000 400128 477012
rect 399536 476972 400128 477000
rect 399536 476960 399542 476972
rect 400122 476960 400128 476972
rect 400180 477000 400186 477012
rect 418154 477000 418160 477012
rect 400180 476972 418160 477000
rect 400180 476960 400186 476972
rect 418154 476960 418160 476972
rect 418212 476960 418218 477012
rect 435726 476960 435732 477012
rect 435784 477000 435790 477012
rect 454034 477000 454040 477012
rect 435784 476972 454040 477000
rect 435784 476960 435790 476972
rect 454034 476960 454040 476972
rect 454092 476960 454098 477012
rect 70210 476892 70216 476944
rect 70268 476932 70274 476944
rect 88702 476932 88708 476944
rect 70268 476904 88708 476932
rect 70268 476892 70274 476904
rect 88702 476892 88708 476904
rect 88760 476932 88766 476944
rect 88760 476904 89714 476932
rect 88760 476892 88766 476904
rect 81802 476864 81808 476876
rect 64846 476836 81808 476864
rect 81802 476824 81808 476836
rect 81860 476864 81866 476876
rect 82630 476864 82636 476876
rect 81860 476836 82636 476864
rect 81860 476824 81866 476836
rect 82630 476824 82636 476836
rect 82688 476824 82694 476876
rect 89686 476864 89714 476904
rect 91094 476892 91100 476944
rect 91152 476932 91158 476944
rect 92198 476932 92204 476944
rect 91152 476904 92204 476932
rect 91152 476892 91158 476904
rect 92198 476892 92204 476904
rect 92256 476932 92262 476944
rect 92256 476904 218744 476932
rect 92256 476892 92262 476904
rect 218716 476876 218744 476904
rect 245930 476892 245936 476944
rect 245988 476932 245994 476944
rect 264974 476932 264980 476944
rect 245988 476904 264980 476932
rect 245988 476892 245994 476904
rect 264974 476892 264980 476904
rect 265032 476892 265038 476944
rect 326982 476892 326988 476944
rect 327040 476932 327046 476944
rect 359642 476932 359648 476944
rect 327040 476904 359648 476932
rect 327040 476892 327046 476904
rect 359642 476892 359648 476904
rect 359700 476892 359706 476944
rect 398834 476892 398840 476944
rect 398892 476932 398898 476944
rect 399570 476932 399576 476944
rect 398892 476904 399576 476932
rect 398892 476892 398898 476904
rect 399570 476892 399576 476904
rect 399628 476932 399634 476944
rect 419534 476932 419540 476944
rect 399628 476904 419540 476932
rect 399628 476892 399634 476904
rect 419534 476892 419540 476904
rect 419592 476892 419598 476944
rect 437474 476892 437480 476944
rect 437532 476932 437538 476944
rect 438118 476932 438124 476944
rect 437532 476904 438124 476932
rect 437532 476892 437538 476904
rect 438118 476892 438124 476904
rect 438176 476932 438182 476944
rect 456794 476932 456800 476944
rect 438176 476904 456800 476932
rect 438176 476892 438182 476904
rect 456794 476892 456800 476904
rect 456852 476892 456858 476944
rect 216398 476864 216404 476876
rect 89686 476836 216404 476864
rect 216398 476824 216404 476836
rect 216456 476824 216462 476876
rect 218698 476824 218704 476876
rect 218756 476864 218762 476876
rect 219250 476864 219256 476876
rect 218756 476836 219256 476864
rect 218756 476824 218762 476836
rect 219250 476824 219256 476836
rect 219308 476864 219314 476876
rect 253382 476864 253388 476876
rect 219308 476836 253388 476864
rect 219308 476824 219314 476836
rect 253382 476824 253388 476836
rect 253440 476864 253446 476876
rect 271874 476864 271880 476876
rect 253440 476836 271880 476864
rect 253440 476824 253446 476836
rect 271874 476824 271880 476836
rect 271932 476824 271938 476876
rect 324222 476824 324228 476876
rect 324280 476864 324286 476876
rect 356974 476864 356980 476876
rect 324280 476836 356980 476864
rect 324280 476824 324286 476836
rect 356974 476824 356980 476836
rect 357032 476824 357038 476876
rect 399754 476824 399760 476876
rect 399812 476864 399818 476876
rect 399812 476836 422294 476864
rect 399812 476824 399818 476836
rect 39666 476756 39672 476808
rect 39724 476796 39730 476808
rect 58158 476796 58164 476808
rect 39724 476768 58164 476796
rect 39724 476756 39730 476768
rect 58158 476756 58164 476768
rect 58216 476756 58222 476808
rect 63494 476756 63500 476808
rect 63552 476796 63558 476808
rect 64230 476796 64236 476808
rect 63552 476768 64236 476796
rect 63552 476756 63558 476768
rect 64230 476756 64236 476768
rect 64288 476796 64294 476808
rect 82814 476796 82820 476808
rect 64288 476768 82820 476796
rect 64288 476756 64294 476768
rect 82814 476756 82820 476768
rect 82872 476796 82878 476808
rect 83918 476796 83924 476808
rect 82872 476768 83924 476796
rect 82872 476756 82878 476768
rect 83918 476756 83924 476768
rect 83976 476756 83982 476808
rect 89714 476756 89720 476808
rect 89772 476796 89778 476808
rect 218054 476796 218060 476808
rect 89772 476768 218060 476796
rect 89772 476756 89778 476768
rect 218054 476756 218060 476768
rect 218112 476796 218118 476808
rect 219342 476796 219348 476808
rect 218112 476768 219348 476796
rect 218112 476756 218118 476768
rect 219342 476756 219348 476768
rect 219400 476756 219406 476808
rect 220722 476756 220728 476808
rect 220780 476796 220786 476808
rect 254486 476796 254492 476808
rect 220780 476768 254492 476796
rect 220780 476756 220786 476768
rect 254486 476756 254492 476768
rect 254544 476796 254550 476808
rect 273254 476796 273260 476808
rect 254544 476768 273260 476796
rect 254544 476756 254550 476768
rect 273254 476756 273260 476768
rect 273312 476756 273318 476808
rect 321462 476756 321468 476808
rect 321520 476796 321526 476808
rect 359366 476796 359372 476808
rect 321520 476768 359372 476796
rect 321520 476756 321526 476768
rect 359366 476756 359372 476768
rect 359424 476756 359430 476808
rect 397178 476756 397184 476808
rect 397236 476796 397242 476808
rect 420914 476796 420920 476808
rect 397236 476768 420920 476796
rect 397236 476756 397242 476768
rect 420914 476756 420920 476768
rect 420972 476756 420978 476808
rect 422266 476796 422294 476836
rect 436830 476824 436836 476876
rect 436888 476864 436894 476876
rect 455414 476864 455420 476876
rect 436888 476836 455420 476864
rect 436888 476824 436894 476836
rect 455414 476824 455420 476836
rect 455472 476824 455478 476876
rect 423122 476796 423128 476808
rect 422266 476768 423128 476796
rect 423122 476756 423128 476768
rect 423180 476796 423186 476808
rect 441614 476796 441620 476808
rect 423180 476768 441620 476796
rect 423180 476756 423186 476768
rect 441614 476756 441620 476768
rect 441672 476756 441678 476808
rect 444190 476756 444196 476808
rect 444248 476796 444254 476808
rect 456886 476796 456892 476808
rect 444248 476768 456892 476796
rect 444248 476756 444254 476768
rect 456886 476756 456892 476768
rect 456944 476756 456950 476808
rect 39850 476688 39856 476740
rect 39908 476728 39914 476740
rect 57882 476728 57888 476740
rect 39908 476700 57888 476728
rect 39908 476688 39914 476700
rect 57882 476688 57888 476700
rect 57940 476688 57946 476740
rect 64874 476688 64880 476740
rect 64932 476728 64938 476740
rect 84010 476728 84016 476740
rect 64932 476700 84016 476728
rect 64932 476688 64938 476700
rect 84010 476688 84016 476700
rect 84068 476688 84074 476740
rect 211706 476688 211712 476740
rect 211764 476728 211770 476740
rect 219158 476728 219164 476740
rect 211764 476700 219164 476728
rect 211764 476688 211770 476700
rect 219158 476688 219164 476700
rect 219216 476728 219222 476740
rect 243170 476728 243176 476740
rect 219216 476700 243176 476728
rect 219216 476688 219222 476700
rect 243170 476688 243176 476700
rect 243228 476728 243234 476740
rect 260834 476728 260840 476740
rect 243228 476700 260840 476728
rect 243228 476688 243234 476700
rect 260834 476688 260840 476700
rect 260892 476688 260898 476740
rect 318702 476688 318708 476740
rect 318760 476728 318766 476740
rect 359550 476728 359556 476740
rect 318760 476700 359556 476728
rect 318760 476688 318766 476700
rect 359550 476688 359556 476700
rect 359608 476688 359614 476740
rect 425514 476688 425520 476740
rect 425572 476728 425578 476740
rect 442994 476728 443000 476740
rect 425572 476700 443000 476728
rect 425572 476688 425578 476700
rect 442994 476688 443000 476700
rect 443052 476688 443058 476740
rect 67542 476620 67548 476672
rect 67600 476660 67606 476672
rect 85298 476660 85304 476672
rect 67600 476632 85304 476660
rect 67600 476620 67606 476632
rect 85298 476620 85304 476632
rect 85356 476660 85362 476672
rect 91278 476660 91284 476672
rect 85356 476632 91284 476660
rect 85356 476620 85362 476632
rect 91278 476620 91284 476632
rect 91336 476620 91342 476672
rect 248598 476660 248604 476672
rect 238726 476632 248604 476660
rect 78214 476552 78220 476604
rect 78272 476592 78278 476604
rect 78272 476564 91232 476592
rect 78272 476552 78278 476564
rect 73154 476484 73160 476536
rect 73212 476524 73218 476536
rect 91094 476524 91100 476536
rect 73212 476496 91100 476524
rect 73212 476484 73218 476496
rect 91094 476484 91100 476496
rect 91152 476484 91158 476536
rect 73798 476416 73804 476468
rect 73856 476456 73862 476468
rect 91204 476456 91232 476564
rect 93026 476484 93032 476536
rect 93084 476524 93090 476536
rect 219802 476524 219808 476536
rect 93084 476496 219808 476524
rect 93084 476484 93090 476496
rect 219802 476484 219808 476496
rect 219860 476524 219866 476536
rect 220722 476524 220728 476536
rect 219860 476496 220728 476524
rect 219860 476484 219866 476496
rect 220722 476484 220728 476496
rect 220780 476484 220786 476536
rect 94406 476456 94412 476468
rect 73856 476428 80054 476456
rect 91204 476428 94412 476456
rect 73856 476416 73862 476428
rect 80026 476252 80054 476428
rect 94406 476416 94412 476428
rect 94464 476456 94470 476468
rect 210602 476456 210608 476468
rect 94464 476428 210608 476456
rect 94464 476416 94470 476428
rect 210602 476416 210608 476428
rect 210660 476456 210666 476468
rect 214558 476456 214564 476468
rect 210660 476428 214564 476456
rect 210660 476416 210666 476428
rect 214558 476416 214564 476428
rect 214616 476416 214622 476468
rect 216490 476416 216496 476468
rect 216548 476456 216554 476468
rect 217042 476456 217048 476468
rect 216548 476428 217048 476456
rect 216548 476416 216554 476428
rect 217042 476416 217048 476428
rect 217100 476456 217106 476468
rect 217100 476428 219434 476456
rect 217100 476416 217106 476428
rect 91186 476348 91192 476400
rect 91244 476388 91250 476400
rect 207014 476388 207020 476400
rect 91244 476360 207020 476388
rect 91244 476348 91250 476360
rect 207014 476348 207020 476360
rect 207072 476348 207078 476400
rect 214374 476348 214380 476400
rect 214432 476388 214438 476400
rect 214432 476360 217824 476388
rect 214432 476348 214438 476360
rect 84010 476280 84016 476332
rect 84068 476320 84074 476332
rect 210786 476320 210792 476332
rect 84068 476292 210792 476320
rect 84068 476280 84074 476292
rect 210786 476280 210792 476292
rect 210844 476320 210850 476332
rect 214834 476320 214840 476332
rect 210844 476292 214840 476320
rect 210844 476280 210850 476292
rect 214834 476280 214840 476292
rect 214892 476280 214898 476332
rect 217796 476264 217824 476360
rect 219406 476320 219434 476428
rect 238726 476320 238754 476632
rect 248598 476620 248604 476632
rect 248656 476660 248662 476672
rect 266354 476660 266360 476672
rect 248656 476632 266360 476660
rect 248656 476620 248662 476632
rect 266354 476620 266360 476632
rect 266412 476620 266418 476672
rect 315942 476620 315948 476672
rect 316000 476660 316006 476672
rect 358170 476660 358176 476672
rect 316000 476632 358176 476660
rect 316000 476620 316006 476632
rect 358170 476620 358176 476632
rect 358228 476620 358234 476672
rect 434438 476620 434444 476672
rect 434496 476660 434502 476672
rect 451366 476660 451372 476672
rect 434496 476632 451372 476660
rect 434496 476620 434502 476632
rect 451366 476620 451372 476632
rect 451424 476620 451430 476672
rect 251082 476552 251088 476604
rect 251140 476592 251146 476604
rect 268194 476592 268200 476604
rect 251140 476564 268200 476592
rect 251140 476552 251146 476564
rect 268194 476552 268200 476564
rect 268252 476552 268258 476604
rect 314562 476552 314568 476604
rect 314620 476592 314626 476604
rect 359458 476592 359464 476604
rect 314620 476564 359464 476592
rect 314620 476552 314626 476564
rect 359458 476552 359464 476564
rect 359516 476552 359522 476604
rect 395798 476552 395804 476604
rect 395856 476592 395862 476604
rect 437474 476592 437480 476604
rect 395856 476564 437480 476592
rect 395856 476552 395862 476564
rect 437474 476552 437480 476564
rect 437532 476552 437538 476604
rect 244274 476484 244280 476536
rect 244332 476524 244338 476536
rect 262214 476524 262220 476536
rect 244332 476496 262220 476524
rect 244332 476484 244338 476496
rect 262214 476484 262220 476496
rect 262272 476484 262278 476536
rect 311802 476484 311808 476536
rect 311860 476524 311866 476536
rect 358078 476524 358084 476536
rect 311860 476496 358084 476524
rect 311860 476484 311866 476496
rect 358078 476484 358084 476496
rect 358136 476484 358142 476536
rect 397822 476484 397828 476536
rect 397880 476524 397886 476536
rect 436830 476524 436836 476536
rect 397880 476496 436836 476524
rect 397880 476484 397886 476496
rect 436830 476484 436836 476496
rect 436888 476484 436894 476536
rect 309042 476416 309048 476468
rect 309100 476456 309106 476468
rect 357158 476456 357164 476468
rect 309100 476428 357164 476456
rect 309100 476416 309106 476428
rect 357158 476416 357164 476428
rect 357216 476416 357222 476468
rect 426158 476416 426164 476468
rect 426216 476456 426222 476468
rect 441982 476456 441988 476468
rect 426216 476428 441988 476456
rect 426216 476416 426222 476428
rect 441982 476416 441988 476428
rect 442040 476416 442046 476468
rect 306098 476348 306104 476400
rect 306156 476388 306162 476400
rect 360194 476388 360200 476400
rect 306156 476360 360200 476388
rect 306156 476348 306162 476360
rect 360194 476348 360200 476360
rect 360252 476348 360258 476400
rect 397730 476348 397736 476400
rect 397788 476388 397794 476400
rect 435726 476388 435732 476400
rect 397788 476360 435732 476388
rect 397788 476348 397794 476360
rect 435726 476348 435732 476360
rect 435784 476348 435790 476400
rect 219406 476292 238754 476320
rect 303522 476280 303528 476332
rect 303580 476320 303586 476332
rect 360286 476320 360292 476332
rect 303580 476292 360292 476320
rect 303580 476280 303586 476292
rect 360286 476280 360292 476292
rect 360344 476280 360350 476332
rect 434622 476280 434628 476332
rect 434680 476320 434686 476332
rect 449894 476320 449900 476332
rect 434680 476292 449900 476320
rect 434680 476280 434686 476292
rect 449894 476280 449900 476292
rect 449952 476280 449958 476332
rect 91186 476252 91192 476264
rect 80026 476224 91192 476252
rect 91186 476212 91192 476224
rect 91244 476212 91250 476264
rect 91278 476212 91284 476264
rect 91336 476252 91342 476264
rect 213454 476252 213460 476264
rect 91336 476224 213460 476252
rect 91336 476212 91342 476224
rect 213454 476212 213460 476224
rect 213512 476252 213518 476264
rect 215110 476252 215116 476264
rect 213512 476224 215116 476252
rect 213512 476212 213518 476224
rect 215110 476212 215116 476224
rect 215168 476212 215174 476264
rect 217778 476212 217784 476264
rect 217836 476252 217842 476264
rect 247126 476252 247132 476264
rect 217836 476224 247132 476252
rect 217836 476212 217842 476224
rect 247126 476212 247132 476224
rect 247184 476212 247190 476264
rect 302142 476212 302148 476264
rect 302200 476252 302206 476264
rect 361666 476252 361672 476264
rect 302200 476224 361672 476252
rect 302200 476212 302206 476224
rect 361666 476212 361672 476224
rect 361724 476212 361730 476264
rect 394050 476212 394056 476264
rect 394108 476252 394114 476264
rect 397730 476252 397736 476264
rect 394108 476224 397736 476252
rect 394108 476212 394114 476224
rect 397730 476212 397736 476224
rect 397788 476212 397794 476264
rect 398926 476212 398932 476264
rect 398984 476252 398990 476264
rect 399662 476252 399668 476264
rect 398984 476224 399668 476252
rect 398984 476212 398990 476224
rect 399662 476212 399668 476224
rect 399720 476212 399726 476264
rect 82630 476144 82636 476196
rect 82688 476184 82694 476196
rect 211706 476184 211712 476196
rect 82688 476156 211712 476184
rect 82688 476144 82694 476156
rect 211706 476144 211712 476156
rect 211764 476144 211770 476196
rect 214742 476144 214748 476196
rect 214800 476184 214806 476196
rect 216398 476184 216404 476196
rect 214800 476156 216404 476184
rect 214800 476144 214806 476156
rect 216398 476144 216404 476156
rect 216456 476184 216462 476196
rect 259362 476184 259368 476196
rect 216456 476156 259368 476184
rect 216456 476144 216462 476156
rect 259362 476144 259368 476156
rect 259420 476144 259426 476196
rect 299382 476144 299388 476196
rect 299440 476184 299446 476196
rect 359274 476184 359280 476196
rect 299440 476156 359280 476184
rect 299440 476144 299446 476156
rect 359274 476144 359280 476156
rect 359332 476144 359338 476196
rect 394142 476144 394148 476196
rect 394200 476184 394206 476196
rect 395798 476184 395804 476196
rect 394200 476156 395804 476184
rect 394200 476144 394206 476156
rect 395798 476144 395804 476156
rect 395856 476144 395862 476196
rect 399202 476144 399208 476196
rect 399260 476184 399266 476196
rect 399846 476184 399852 476196
rect 399260 476156 399852 476184
rect 399260 476144 399266 476156
rect 399846 476144 399852 476156
rect 399904 476144 399910 476196
rect 83918 476076 83924 476128
rect 83976 476116 83982 476128
rect 217962 476116 217968 476128
rect 83976 476088 217968 476116
rect 83976 476076 83982 476088
rect 217962 476076 217968 476088
rect 218020 476076 218026 476128
rect 296254 476076 296260 476128
rect 296312 476116 296318 476128
rect 357986 476116 357992 476128
rect 296312 476088 357992 476116
rect 296312 476076 296318 476088
rect 357986 476076 357992 476088
rect 358044 476076 358050 476128
rect 394234 476076 394240 476128
rect 394292 476116 394298 476128
rect 397822 476116 397828 476128
rect 394292 476088 397828 476116
rect 394292 476076 394298 476088
rect 397822 476076 397828 476088
rect 397880 476076 397886 476128
rect 399294 476076 399300 476128
rect 399352 476116 399358 476128
rect 399754 476116 399760 476128
rect 399352 476088 399760 476116
rect 399352 476076 399358 476088
rect 399754 476076 399760 476088
rect 399812 476076 399818 476128
rect 400122 476076 400128 476128
rect 400180 476116 400186 476128
rect 433334 476116 433340 476128
rect 400180 476088 433340 476116
rect 400180 476076 400186 476088
rect 433334 476076 433340 476088
rect 433392 476076 433398 476128
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 7558 474756 7564 474768
rect 3108 474728 7564 474756
rect 3108 474716 3114 474728
rect 7558 474716 7564 474728
rect 7616 474716 7622 474768
rect 215846 474648 215852 474700
rect 215904 474688 215910 474700
rect 268010 474688 268016 474700
rect 215904 474660 268016 474688
rect 215904 474648 215910 474660
rect 268010 474648 268016 474660
rect 268068 474648 268074 474700
rect 393958 474648 393964 474700
rect 394016 474688 394022 474700
rect 395062 474688 395068 474700
rect 394016 474660 395068 474688
rect 394016 474648 394022 474660
rect 395062 474648 395068 474660
rect 395120 474648 395126 474700
rect 395430 474648 395436 474700
rect 395488 474688 395494 474700
rect 477494 474688 477500 474700
rect 395488 474660 477500 474688
rect 395488 474648 395494 474660
rect 477494 474648 477500 474660
rect 477552 474648 477558 474700
rect 219066 474580 219072 474632
rect 219124 474620 219130 474632
rect 273254 474620 273260 474632
rect 219124 474592 273260 474620
rect 219124 474580 219130 474592
rect 273254 474580 273260 474592
rect 273312 474580 273318 474632
rect 395614 474580 395620 474632
rect 395672 474620 395678 474632
rect 480530 474620 480536 474632
rect 395672 474592 480536 474620
rect 395672 474580 395678 474592
rect 480530 474580 480536 474592
rect 480588 474580 480594 474632
rect 215938 474512 215944 474564
rect 215996 474552 216002 474564
rect 270494 474552 270500 474564
rect 215996 474524 270500 474552
rect 215996 474512 216002 474524
rect 270494 474512 270500 474524
rect 270552 474512 270558 474564
rect 395706 474512 395712 474564
rect 395764 474552 395770 474564
rect 483014 474552 483020 474564
rect 395764 474524 483020 474552
rect 395764 474512 395770 474524
rect 483014 474512 483020 474524
rect 483072 474512 483078 474564
rect 219710 474444 219716 474496
rect 219768 474484 219774 474496
rect 276014 474484 276020 474496
rect 219768 474456 276020 474484
rect 219768 474444 219774 474456
rect 276014 474444 276020 474456
rect 276072 474444 276078 474496
rect 395798 474444 395804 474496
rect 395856 474484 395862 474496
rect 485774 474484 485780 474496
rect 395856 474456 485780 474484
rect 395856 474444 395862 474456
rect 485774 474444 485780 474456
rect 485832 474444 485838 474496
rect 214834 474376 214840 474428
rect 214892 474416 214898 474428
rect 277578 474416 277584 474428
rect 214892 474388 277584 474416
rect 214892 474376 214898 474388
rect 277578 474376 277584 474388
rect 277636 474376 277642 474428
rect 395982 474376 395988 474428
rect 396040 474416 396046 474428
rect 488534 474416 488540 474428
rect 396040 474388 488540 474416
rect 396040 474376 396046 474388
rect 488534 474376 488540 474388
rect 488592 474376 488598 474428
rect 219618 474308 219624 474360
rect 219676 474348 219682 474360
rect 285674 474348 285680 474360
rect 219676 474320 285680 474348
rect 219676 474308 219682 474320
rect 285674 474308 285680 474320
rect 285732 474308 285738 474360
rect 395890 474308 395896 474360
rect 395948 474348 395954 474360
rect 490466 474348 490472 474360
rect 395948 474320 490472 474348
rect 395948 474308 395954 474320
rect 490466 474308 490472 474320
rect 490524 474308 490530 474360
rect 213086 474240 213092 474292
rect 213144 474280 213150 474292
rect 280154 474280 280160 474292
rect 213144 474252 280160 474280
rect 213144 474240 213150 474252
rect 280154 474240 280160 474252
rect 280212 474240 280218 474292
rect 395246 474240 395252 474292
rect 395304 474280 395310 474292
rect 492674 474280 492680 474292
rect 395304 474252 492680 474280
rect 395304 474240 395310 474252
rect 492674 474240 492680 474252
rect 492732 474240 492738 474292
rect 215754 474172 215760 474224
rect 215812 474212 215818 474224
rect 282914 474212 282920 474224
rect 215812 474184 282920 474212
rect 215812 474172 215818 474184
rect 282914 474172 282920 474184
rect 282972 474172 282978 474224
rect 399478 474172 399484 474224
rect 399536 474212 399542 474224
rect 502334 474212 502340 474224
rect 399536 474184 502340 474212
rect 399536 474172 399542 474184
rect 502334 474172 502340 474184
rect 502392 474172 502398 474224
rect 218698 474104 218704 474156
rect 218756 474144 218762 474156
rect 292574 474144 292580 474156
rect 218756 474116 292580 474144
rect 218756 474104 218762 474116
rect 292574 474104 292580 474116
rect 292632 474104 292638 474156
rect 392394 474104 392400 474156
rect 392452 474144 392458 474156
rect 495434 474144 495440 474156
rect 392452 474116 495440 474144
rect 392452 474104 392458 474116
rect 495434 474104 495440 474116
rect 495492 474104 495498 474156
rect 208946 474036 208952 474088
rect 209004 474076 209010 474088
rect 287698 474076 287704 474088
rect 209004 474048 287704 474076
rect 209004 474036 209010 474048
rect 287698 474036 287704 474048
rect 287756 474036 287762 474088
rect 393038 474036 393044 474088
rect 393096 474076 393102 474088
rect 498194 474076 498200 474088
rect 393096 474048 498200 474076
rect 393096 474036 393102 474048
rect 498194 474036 498200 474048
rect 498252 474036 498258 474088
rect 210326 473968 210332 474020
rect 210384 474008 210390 474020
rect 289814 474008 289820 474020
rect 210384 473980 289820 474008
rect 210384 473968 210390 473980
rect 289814 473968 289820 473980
rect 289872 473968 289878 474020
rect 392946 473968 392952 474020
rect 393004 474008 393010 474020
rect 500954 474008 500960 474020
rect 393004 473980 500960 474008
rect 393004 473968 393010 473980
rect 500954 473968 500960 473980
rect 501012 473968 501018 474020
rect 216030 473900 216036 473952
rect 216088 473940 216094 473952
rect 264974 473940 264980 473952
rect 216088 473912 264980 473940
rect 216088 473900 216094 473912
rect 264974 473900 264980 473912
rect 265032 473900 265038 473952
rect 395522 473900 395528 473952
rect 395580 473940 395586 473952
rect 474734 473940 474740 473952
rect 395580 473912 474740 473940
rect 395580 473900 395586 473912
rect 474734 473900 474740 473912
rect 474792 473900 474798 473952
rect 216214 473832 216220 473884
rect 216272 473872 216278 473884
rect 263594 473872 263600 473884
rect 216272 473844 263600 473872
rect 216272 473832 216278 473844
rect 263594 473832 263600 473844
rect 263652 473832 263658 473884
rect 397914 473832 397920 473884
rect 397972 473872 397978 473884
rect 465074 473872 465080 473884
rect 397972 473844 465080 473872
rect 397972 473832 397978 473844
rect 465074 473832 465080 473844
rect 465132 473832 465138 473884
rect 216306 473764 216312 473816
rect 216364 473804 216370 473816
rect 260834 473804 260840 473816
rect 216364 473776 260840 473804
rect 216364 473764 216370 473776
rect 260834 473764 260840 473776
rect 260892 473764 260898 473816
rect 395062 473764 395068 473816
rect 395120 473804 395126 473816
rect 438854 473804 438860 473816
rect 395120 473776 438860 473804
rect 395120 473764 395126 473776
rect 438854 473764 438860 473776
rect 438912 473764 438918 473816
rect 395154 471928 395160 471980
rect 395212 471968 395218 471980
rect 440234 471968 440240 471980
rect 395212 471940 440240 471968
rect 395212 471928 395218 471940
rect 440234 471928 440240 471940
rect 440292 471928 440298 471980
rect 392486 471452 392492 471504
rect 392544 471492 392550 471504
rect 445754 471492 445760 471504
rect 392544 471464 445760 471492
rect 392544 471452 392550 471464
rect 445754 471452 445760 471464
rect 445812 471452 445818 471504
rect 393222 471384 393228 471436
rect 393280 471424 393286 471436
rect 447134 471424 447140 471436
rect 393280 471396 447140 471424
rect 393280 471384 393286 471396
rect 447134 471384 447140 471396
rect 447192 471384 447198 471436
rect 392762 471316 392768 471368
rect 392820 471356 392826 471368
rect 449894 471356 449900 471368
rect 392820 471328 449900 471356
rect 392820 471316 392826 471328
rect 449894 471316 449900 471328
rect 449952 471316 449958 471368
rect 393130 471248 393136 471300
rect 393188 471288 393194 471300
rect 505094 471288 505100 471300
rect 393188 471260 505100 471288
rect 393188 471248 393194 471260
rect 505094 471248 505100 471260
rect 505152 471248 505158 471300
rect 393866 471180 393872 471232
rect 393924 471220 393930 471232
rect 395154 471220 395160 471232
rect 393924 471192 395160 471220
rect 393924 471180 393930 471192
rect 395154 471180 395160 471192
rect 395212 471180 395218 471232
rect 182910 470568 182916 470620
rect 182968 470608 182974 470620
rect 580166 470608 580172 470620
rect 182968 470580 580172 470608
rect 182968 470568 182974 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 15838 462380 15844 462392
rect 3568 462352 15844 462380
rect 3568 462340 3574 462352
rect 15838 462340 15844 462352
rect 15896 462340 15902 462392
rect 188430 456764 188436 456816
rect 188488 456804 188494 456816
rect 580166 456804 580172 456816
rect 188488 456776 580172 456804
rect 188488 456764 188494 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 358814 454724 358820 454776
rect 358872 454764 358878 454776
rect 359734 454764 359740 454776
rect 358872 454736 359740 454764
rect 358872 454724 358878 454736
rect 359734 454724 359740 454736
rect 359792 454764 359798 454776
rect 538214 454764 538220 454776
rect 359792 454736 538220 454764
rect 359792 454724 359798 454736
rect 538214 454724 538220 454736
rect 538272 454724 538278 454776
rect 216766 454656 216772 454708
rect 216824 454696 216830 454708
rect 217686 454696 217692 454708
rect 216824 454668 217692 454696
rect 216824 454656 216830 454668
rect 217686 454656 217692 454668
rect 217744 454696 217750 454708
rect 396442 454696 396448 454708
rect 217744 454668 396448 454696
rect 217744 454656 217750 454668
rect 396442 454656 396448 454668
rect 396500 454696 396506 454708
rect 396626 454696 396632 454708
rect 396500 454668 396632 454696
rect 396500 454656 396506 454668
rect 396626 454656 396632 454668
rect 396684 454656 396690 454708
rect 179046 453296 179052 453348
rect 179104 453336 179110 453348
rect 358814 453336 358820 453348
rect 179104 453308 358820 453336
rect 179104 453296 179110 453308
rect 358814 453296 358820 453308
rect 358872 453296 358878 453348
rect 214558 451868 214564 451920
rect 214616 451908 214622 451920
rect 249794 451908 249800 451920
rect 214616 451880 249800 451908
rect 214616 451868 214622 451880
rect 249794 451868 249800 451880
rect 249852 451868 249858 451920
rect 216950 450780 216956 450832
rect 217008 450820 217014 450832
rect 217318 450820 217324 450832
rect 217008 450792 217324 450820
rect 217008 450780 217014 450792
rect 217318 450780 217324 450792
rect 217376 450780 217382 450832
rect 217318 450508 217324 450560
rect 217376 450548 217382 450560
rect 396534 450548 396540 450560
rect 217376 450520 396540 450548
rect 217376 450508 217382 450520
rect 396534 450508 396540 450520
rect 396592 450508 396598 450560
rect 210142 449216 210148 449268
rect 210200 449256 210206 449268
rect 247034 449256 247040 449268
rect 210200 449228 247040 449256
rect 210200 449216 210206 449228
rect 247034 449216 247040 449228
rect 247092 449216 247098 449268
rect 71682 449148 71688 449200
rect 71740 449188 71746 449200
rect 212534 449188 212540 449200
rect 71740 449160 212540 449188
rect 71740 449148 71746 449160
rect 212534 449148 212540 449160
rect 212592 449148 212598 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 14550 448576 14556 448588
rect 3200 448548 14556 448576
rect 3200 448536 3206 448548
rect 14550 448536 14556 448548
rect 14608 448536 14614 448588
rect 142062 448468 142068 448520
rect 142120 448508 142126 448520
rect 209222 448508 209228 448520
rect 142120 448480 209228 448508
rect 142120 448468 142126 448480
rect 209222 448468 209228 448480
rect 209280 448468 209286 448520
rect 139302 448400 139308 448452
rect 139360 448440 139366 448452
rect 209406 448440 209412 448452
rect 139360 448412 209412 448440
rect 139360 448400 139366 448412
rect 209406 448400 209412 448412
rect 209464 448400 209470 448452
rect 136542 448332 136548 448384
rect 136600 448372 136606 448384
rect 209038 448372 209044 448384
rect 136600 448344 209044 448372
rect 136600 448332 136606 448344
rect 209038 448332 209044 448344
rect 209096 448332 209102 448384
rect 133782 448264 133788 448316
rect 133840 448304 133846 448316
rect 209590 448304 209596 448316
rect 133840 448276 209596 448304
rect 133840 448264 133846 448276
rect 209590 448264 209596 448276
rect 209648 448264 209654 448316
rect 131022 448196 131028 448248
rect 131080 448236 131086 448248
rect 209498 448236 209504 448248
rect 131080 448208 209504 448236
rect 131080 448196 131086 448208
rect 209498 448196 209504 448208
rect 209556 448196 209562 448248
rect 91002 448128 91008 448180
rect 91060 448168 91066 448180
rect 206554 448168 206560 448180
rect 91060 448140 206560 448168
rect 91060 448128 91066 448140
rect 206554 448128 206560 448140
rect 206612 448128 206618 448180
rect 88242 448060 88248 448112
rect 88300 448100 88306 448112
rect 206646 448100 206652 448112
rect 88300 448072 206652 448100
rect 88300 448060 88306 448072
rect 206646 448060 206652 448072
rect 206704 448060 206710 448112
rect 86862 447992 86868 448044
rect 86920 448032 86926 448044
rect 206738 448032 206744 448044
rect 86920 448004 206744 448032
rect 86920 447992 86926 448004
rect 206738 447992 206744 448004
rect 206796 447992 206802 448044
rect 84102 447924 84108 447976
rect 84160 447964 84166 447976
rect 206462 447964 206468 447976
rect 84160 447936 206468 447964
rect 84160 447924 84166 447936
rect 206462 447924 206468 447936
rect 206520 447924 206526 447976
rect 81342 447856 81348 447908
rect 81400 447896 81406 447908
rect 206370 447896 206376 447908
rect 81400 447868 206376 447896
rect 81400 447856 81406 447868
rect 206370 447856 206376 447868
rect 206428 447856 206434 447908
rect 78582 447788 78588 447840
rect 78640 447828 78646 447840
rect 206278 447828 206284 447840
rect 78640 447800 206284 447828
rect 78640 447788 78646 447800
rect 206278 447788 206284 447800
rect 206336 447788 206342 447840
rect 143442 447720 143448 447772
rect 143500 447760 143506 447772
rect 209314 447760 209320 447772
rect 143500 447732 209320 447760
rect 143500 447720 143506 447732
rect 209314 447720 209320 447732
rect 209372 447720 209378 447772
rect 146202 447652 146208 447704
rect 146260 447692 146266 447704
rect 209130 447692 209136 447704
rect 146260 447664 209136 447692
rect 146260 447652 146266 447664
rect 209130 447652 209136 447664
rect 209188 447652 209194 447704
rect 170858 447040 170864 447092
rect 170916 447080 170922 447092
rect 180150 447080 180156 447092
rect 170916 447052 180156 447080
rect 170916 447040 170922 447052
rect 180150 447040 180156 447052
rect 180208 447040 180214 447092
rect 351086 447040 351092 447092
rect 351144 447080 351150 447092
rect 374638 447080 374644 447092
rect 351144 447052 374644 447080
rect 351144 447040 351150 447052
rect 374638 447040 374644 447052
rect 374696 447040 374702 447092
rect 530486 446972 530492 447024
rect 530544 447012 530550 447024
rect 536834 447012 536840 447024
rect 530544 446984 536840 447012
rect 530544 446972 530550 446984
rect 536834 446972 536840 446984
rect 536892 446972 536898 447024
rect 218974 446360 218980 446412
rect 219032 446400 219038 446412
rect 252554 446400 252560 446412
rect 219032 446372 252560 446400
rect 219032 446360 219038 446372
rect 252554 446360 252560 446372
rect 252612 446360 252618 446412
rect 124122 445680 124128 445732
rect 124180 445720 124186 445732
rect 212258 445720 212264 445732
rect 124180 445692 212264 445720
rect 124180 445680 124186 445692
rect 212258 445680 212264 445692
rect 212316 445680 212322 445732
rect 121362 445612 121368 445664
rect 121420 445652 121426 445664
rect 212166 445652 212172 445664
rect 121420 445624 212172 445652
rect 121420 445612 121426 445624
rect 212166 445612 212172 445624
rect 212224 445612 212230 445664
rect 118602 445544 118608 445596
rect 118660 445584 118666 445596
rect 211982 445584 211988 445596
rect 118660 445556 211988 445584
rect 118660 445544 118666 445556
rect 211982 445544 211988 445556
rect 212040 445544 212046 445596
rect 117222 445476 117228 445528
rect 117280 445516 117286 445528
rect 211798 445516 211804 445528
rect 117280 445488 211804 445516
rect 117280 445476 117286 445488
rect 211798 445476 211804 445488
rect 211856 445476 211862 445528
rect 114462 445408 114468 445460
rect 114520 445448 114526 445460
rect 211890 445448 211896 445460
rect 114520 445420 211896 445448
rect 114520 445408 114526 445420
rect 211890 445408 211896 445420
rect 211948 445408 211954 445460
rect 106182 445340 106188 445392
rect 106240 445380 106246 445392
rect 215018 445380 215024 445392
rect 106240 445352 215024 445380
rect 106240 445340 106246 445352
rect 215018 445340 215024 445352
rect 215076 445340 215082 445392
rect 104802 445272 104808 445324
rect 104860 445312 104866 445324
rect 214466 445312 214472 445324
rect 104860 445284 214472 445312
rect 104860 445272 104866 445284
rect 214466 445272 214472 445284
rect 214524 445272 214530 445324
rect 102042 445204 102048 445256
rect 102100 445244 102106 445256
rect 214282 445244 214288 445256
rect 102100 445216 214288 445244
rect 102100 445204 102106 445216
rect 214282 445204 214288 445216
rect 214340 445204 214346 445256
rect 99282 445136 99288 445188
rect 99340 445176 99346 445188
rect 214742 445176 214748 445188
rect 99340 445148 214748 445176
rect 99340 445136 99346 445148
rect 214742 445136 214748 445148
rect 214800 445136 214806 445188
rect 96522 445068 96528 445120
rect 96580 445108 96586 445120
rect 214650 445108 214656 445120
rect 96580 445080 214656 445108
rect 96580 445068 96586 445080
rect 214650 445068 214656 445080
rect 214708 445068 214714 445120
rect 68922 445000 68928 445052
rect 68980 445040 68986 445052
rect 208578 445040 208584 445052
rect 68980 445012 208584 445040
rect 68980 445000 68986 445012
rect 208578 445000 208584 445012
rect 208636 445000 208642 445052
rect 126882 444932 126888 444984
rect 126940 444972 126946 444984
rect 212074 444972 212080 444984
rect 126940 444944 212080 444972
rect 126940 444932 126946 444944
rect 212074 444932 212080 444944
rect 212132 444932 212138 444984
rect 129642 444864 129648 444916
rect 129700 444904 129706 444916
rect 209682 444904 209688 444916
rect 129700 444876 209688 444904
rect 129700 444864 129706 444876
rect 209682 444864 209688 444876
rect 209740 444864 209746 444916
rect 178494 444320 178500 444372
rect 178552 444360 178558 444372
rect 179046 444360 179052 444372
rect 178552 444332 179052 444360
rect 178552 444320 178558 444332
rect 179046 444320 179052 444332
rect 179104 444320 179110 444372
rect 77202 443640 77208 443692
rect 77260 443680 77266 443692
rect 219894 443680 219900 443692
rect 77260 443652 219900 443680
rect 77260 443640 77266 443652
rect 219894 443640 219900 443652
rect 219952 443640 219958 443692
rect 38470 443232 38476 443284
rect 38528 443272 38534 443284
rect 178494 443272 178500 443284
rect 38528 443244 178500 443272
rect 38528 443232 38534 443244
rect 178494 443232 178500 443244
rect 178552 443232 178558 443284
rect 548518 430584 548524 430636
rect 548576 430624 548582 430636
rect 580166 430624 580172 430636
rect 548576 430596 580172 430624
rect 548576 430584 548582 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 10318 422328 10324 422340
rect 3568 422300 10324 422328
rect 3568 422288 3574 422300
rect 10318 422288 10324 422300
rect 10376 422288 10382 422340
rect 540330 404336 540336 404388
rect 540388 404376 540394 404388
rect 580166 404376 580172 404388
rect 540388 404348 580172 404376
rect 540388 404336 540394 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 11790 397508 11796 397520
rect 3384 397480 11796 397508
rect 3384 397468 3390 397480
rect 11790 397468 11796 397480
rect 11848 397468 11854 397520
rect 217594 393320 217600 393372
rect 217652 393360 217658 393372
rect 218054 393360 218060 393372
rect 217652 393332 218060 393360
rect 217652 393320 217658 393332
rect 218054 393320 218060 393332
rect 218112 393320 218118 393372
rect 217318 392028 217324 392080
rect 217376 392068 217382 392080
rect 218698 392068 218704 392080
rect 217376 392040 218704 392068
rect 217376 392028 217382 392040
rect 218698 392028 218704 392040
rect 218756 392028 218762 392080
rect 218514 391960 218520 392012
rect 218572 392000 218578 392012
rect 218572 391972 218744 392000
rect 218572 391960 218578 391972
rect 218716 391944 218744 391972
rect 218698 391892 218704 391944
rect 218756 391892 218762 391944
rect 547138 378156 547144 378208
rect 547196 378196 547202 378208
rect 580166 378196 580172 378208
rect 547196 378168 580172 378196
rect 547196 378156 547202 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 10410 371260 10416 371272
rect 3384 371232 10416 371260
rect 3384 371220 3390 371232
rect 10410 371220 10416 371232
rect 10468 371220 10474 371272
rect 362218 367140 362224 367192
rect 362276 367180 362282 367192
rect 396718 367180 396724 367192
rect 362276 367152 396724 367180
rect 362276 367140 362282 367152
rect 396718 367140 396724 367152
rect 396776 367140 396782 367192
rect 358262 367072 358268 367124
rect 358320 367112 358326 367124
rect 396534 367112 396540 367124
rect 358320 367084 396540 367112
rect 358320 367072 358326 367084
rect 396534 367072 396540 367084
rect 396592 367072 396598 367124
rect 396442 367004 396448 367056
rect 396500 367044 396506 367056
rect 396718 367044 396724 367056
rect 396500 367016 396724 367044
rect 396500 367004 396506 367016
rect 396718 367004 396724 367016
rect 396776 367004 396782 367056
rect 542998 364352 543004 364404
rect 543056 364392 543062 364404
rect 579798 364392 579804 364404
rect 543056 364364 579804 364392
rect 543056 364352 543062 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 38194 360000 38200 360052
rect 38252 360040 38258 360052
rect 38252 360012 200114 360040
rect 38252 360000 38258 360012
rect 200086 359972 200114 360012
rect 218606 360000 218612 360052
rect 218664 360040 218670 360052
rect 224218 360040 224224 360052
rect 218664 360012 224224 360040
rect 218664 360000 218670 360012
rect 224218 360000 224224 360012
rect 224276 360000 224282 360052
rect 234062 360000 234068 360052
rect 234120 360040 234126 360052
rect 396626 360040 396632 360052
rect 234120 360012 396632 360040
rect 234120 360000 234126 360012
rect 396626 360000 396632 360012
rect 396684 360000 396690 360052
rect 218514 359972 218520 359984
rect 200086 359944 218520 359972
rect 218514 359932 218520 359944
rect 218572 359972 218578 359984
rect 218572 359944 361620 359972
rect 218572 359932 218578 359944
rect 210970 359864 210976 359916
rect 211028 359904 211034 359916
rect 270494 359904 270500 359916
rect 211028 359876 270500 359904
rect 211028 359864 211034 359876
rect 270494 359864 270500 359876
rect 270552 359864 270558 359916
rect 311710 359864 311716 359916
rect 311768 359904 311774 359916
rect 357894 359904 357900 359916
rect 311768 359876 357900 359904
rect 311768 359864 311774 359876
rect 357894 359864 357900 359876
rect 357952 359864 357958 359916
rect 361592 359848 361620 359944
rect 212442 359796 212448 359848
rect 212500 359836 212506 359848
rect 273438 359836 273444 359848
rect 212500 359808 273444 359836
rect 212500 359796 212506 359808
rect 273438 359796 273444 359808
rect 273496 359796 273502 359848
rect 279326 359796 279332 359848
rect 279384 359836 279390 359848
rect 357802 359836 357808 359848
rect 279384 359808 357808 359836
rect 279384 359796 279390 359808
rect 357802 359796 357808 359808
rect 357860 359796 357866 359848
rect 361574 359796 361580 359848
rect 361632 359836 361638 359848
rect 362218 359836 362224 359848
rect 361632 359808 362224 359836
rect 361632 359796 361638 359808
rect 362218 359796 362224 359808
rect 362276 359796 362282 359848
rect 393774 359796 393780 359848
rect 393832 359836 393838 359848
rect 394142 359836 394148 359848
rect 393832 359808 394148 359836
rect 393832 359796 393838 359808
rect 394142 359796 394148 359808
rect 394200 359796 394206 359848
rect 215202 359728 215208 359780
rect 215260 359768 215266 359780
rect 276382 359768 276388 359780
rect 215260 359740 276388 359768
rect 215260 359728 215266 359740
rect 276382 359728 276388 359740
rect 276440 359728 276446 359780
rect 300670 359728 300676 359780
rect 300728 359768 300734 359780
rect 395246 359768 395252 359780
rect 300728 359740 395252 359768
rect 300728 359728 300734 359740
rect 395246 359728 395252 359740
rect 395304 359728 395310 359780
rect 210326 359660 210332 359712
rect 210384 359700 210390 359712
rect 273070 359700 273076 359712
rect 210384 359672 273076 359700
rect 210384 359660 210390 359672
rect 273070 359660 273076 359672
rect 273128 359660 273134 359712
rect 277118 359660 277124 359712
rect 277176 359700 277182 359712
rect 398006 359700 398012 359712
rect 277176 359672 398012 359700
rect 277176 359660 277182 359672
rect 398006 359660 398012 359672
rect 398064 359660 398070 359712
rect 208946 359592 208952 359644
rect 209004 359632 209010 359644
rect 270126 359632 270132 359644
rect 209004 359604 270132 359632
rect 209004 359592 209010 359604
rect 270126 359592 270132 359604
rect 270184 359592 270190 359644
rect 271230 359592 271236 359644
rect 271288 359632 271294 359644
rect 397822 359632 397828 359644
rect 271288 359604 397828 359632
rect 271288 359592 271294 359604
rect 397822 359592 397828 359604
rect 397880 359592 397886 359644
rect 215754 359524 215760 359576
rect 215812 359564 215818 359576
rect 263502 359564 263508 359576
rect 215812 359536 263508 359564
rect 215812 359524 215818 359536
rect 263502 359524 263508 359536
rect 263560 359524 263566 359576
rect 264606 359524 264612 359576
rect 264664 359564 264670 359576
rect 398190 359564 398196 359576
rect 264664 359536 398196 359564
rect 264664 359524 264670 359536
rect 398190 359524 398196 359536
rect 398248 359524 398254 359576
rect 213086 359456 213092 359508
rect 213144 359496 213150 359508
rect 259730 359496 259736 359508
rect 213144 359468 259736 359496
rect 213144 359456 213150 359468
rect 259730 359456 259736 359468
rect 259788 359456 259794 359508
rect 261294 359456 261300 359508
rect 261352 359496 261358 359508
rect 398558 359496 398564 359508
rect 261352 359468 398564 359496
rect 261352 359456 261358 359468
rect 398558 359456 398564 359468
rect 398616 359456 398622 359508
rect 217318 359388 217324 359440
rect 217376 359428 217382 359440
rect 276106 359428 276112 359440
rect 217376 359400 276112 359428
rect 217376 359388 217382 359400
rect 276106 359388 276112 359400
rect 276164 359388 276170 359440
rect 314286 359388 314292 359440
rect 314344 359428 314350 359440
rect 359642 359428 359648 359440
rect 314344 359400 359648 359428
rect 314344 359388 314350 359400
rect 359642 359388 359648 359400
rect 359700 359388 359706 359440
rect 219618 359320 219624 359372
rect 219676 359360 219682 359372
rect 266814 359360 266820 359372
rect 219676 359332 266820 359360
rect 219676 359320 219682 359332
rect 266814 359320 266820 359332
rect 266872 359320 266878 359372
rect 397362 359320 397368 359372
rect 397420 359320 397426 359372
rect 211062 359252 211068 359304
rect 211120 359292 211126 359304
rect 257246 359292 257252 359304
rect 211120 359264 257252 359292
rect 211120 359252 211126 359264
rect 257246 359252 257252 359264
rect 257304 359252 257310 359304
rect 214834 359184 214840 359236
rect 214892 359224 214898 359236
rect 256878 359224 256884 359236
rect 214892 359196 256884 359224
rect 214892 359184 214898 359196
rect 256878 359184 256884 359196
rect 256936 359184 256942 359236
rect 397270 359116 397276 359168
rect 397328 359156 397334 359168
rect 397380 359156 397408 359320
rect 397328 359128 397408 359156
rect 397328 359116 397334 359128
rect 217226 358708 217232 358760
rect 217284 358748 217290 358760
rect 396810 358748 396816 358760
rect 217284 358720 396816 358748
rect 217284 358708 217290 358720
rect 396810 358708 396816 358720
rect 396868 358708 396874 358760
rect 216950 358640 216956 358692
rect 217008 358680 217014 358692
rect 217318 358680 217324 358692
rect 217008 358652 217324 358680
rect 217008 358640 217014 358652
rect 217318 358640 217324 358652
rect 217376 358680 217382 358692
rect 397086 358680 397092 358692
rect 217376 358652 397092 358680
rect 217376 358640 217382 358652
rect 397086 358640 397092 358652
rect 397144 358640 397150 358692
rect 217870 358572 217876 358624
rect 217928 358612 217934 358624
rect 396902 358612 396908 358624
rect 217928 358584 396908 358612
rect 217928 358572 217934 358584
rect 396902 358572 396908 358584
rect 396960 358572 396966 358624
rect 218330 358504 218336 358556
rect 218388 358544 218394 358556
rect 235994 358544 236000 358556
rect 218388 358516 236000 358544
rect 218388 358504 218394 358516
rect 235994 358504 236000 358516
rect 236052 358504 236058 358556
rect 305454 358504 305460 358556
rect 305512 358544 305518 358556
rect 359550 358544 359556 358556
rect 305512 358516 359556 358544
rect 305512 358504 305518 358516
rect 359550 358504 359556 358516
rect 359608 358504 359614 358556
rect 216030 358436 216036 358488
rect 216088 358476 216094 358488
rect 239950 358476 239956 358488
rect 216088 358448 239956 358476
rect 216088 358436 216094 358448
rect 239950 358436 239956 358448
rect 240008 358436 240014 358488
rect 302510 358436 302516 358488
rect 302568 358476 302574 358488
rect 358170 358476 358176 358488
rect 302568 358448 358176 358476
rect 302568 358436 302574 358448
rect 358170 358436 358176 358448
rect 358228 358436 358234 358488
rect 215846 358368 215852 358420
rect 215904 358408 215910 358420
rect 243630 358408 243636 358420
rect 215904 358380 243636 358408
rect 215904 358368 215910 358380
rect 243630 358368 243636 358380
rect 243688 358368 243694 358420
rect 302878 358368 302884 358420
rect 302936 358408 302942 358420
rect 359182 358408 359188 358420
rect 302936 358380 359188 358408
rect 302936 358368 302942 358380
rect 359182 358368 359188 358380
rect 359240 358368 359246 358420
rect 215938 358300 215944 358352
rect 215996 358340 216002 358352
rect 246942 358340 246948 358352
rect 215996 358312 246948 358340
rect 215996 358300 216002 358312
rect 246942 358300 246948 358312
rect 247000 358300 247006 358352
rect 299566 358300 299572 358352
rect 299624 358340 299630 358352
rect 359458 358340 359464 358352
rect 299624 358312 359464 358340
rect 299624 358300 299630 358312
rect 359458 358300 359464 358312
rect 359516 358300 359522 358352
rect 147582 358232 147588 358284
rect 147640 358272 147646 358284
rect 178402 358272 178408 358284
rect 147640 358244 178408 358272
rect 147640 358232 147646 358244
rect 178402 358232 178408 358244
rect 178460 358232 178466 358284
rect 219066 358232 219072 358284
rect 219124 358272 219130 358284
rect 250254 358272 250260 358284
rect 219124 358244 250260 358272
rect 219124 358232 219130 358244
rect 250254 358232 250260 358244
rect 250312 358232 250318 358284
rect 296622 358232 296628 358284
rect 296680 358272 296686 358284
rect 358078 358272 358084 358284
rect 296680 358244 358084 358272
rect 296680 358232 296686 358244
rect 358078 358232 358084 358244
rect 358136 358232 358142 358284
rect 146846 358164 146852 358216
rect 146904 358204 146910 358216
rect 178310 358204 178316 358216
rect 146904 358176 178316 358204
rect 146904 358164 146910 358176
rect 178310 358164 178316 358176
rect 178368 358164 178374 358216
rect 219710 358164 219716 358216
rect 219768 358204 219774 358216
rect 253566 358204 253572 358216
rect 219768 358176 253572 358204
rect 219768 358164 219774 358176
rect 253566 358164 253572 358176
rect 253624 358164 253630 358216
rect 293678 358164 293684 358216
rect 293736 358204 293742 358216
rect 357158 358204 357164 358216
rect 293736 358176 357164 358204
rect 293736 358164 293742 358176
rect 357158 358164 357164 358176
rect 357216 358164 357222 358216
rect 146478 358096 146484 358148
rect 146536 358136 146542 358148
rect 186958 358136 186964 358148
rect 146536 358108 186964 358136
rect 146536 358096 146542 358108
rect 186958 358096 186964 358108
rect 187016 358096 187022 358148
rect 216214 358096 216220 358148
rect 216272 358136 216278 358148
rect 235902 358136 235908 358148
rect 216272 358108 235908 358136
rect 216272 358096 216278 358108
rect 235902 358096 235908 358108
rect 235960 358096 235966 358148
rect 235994 358096 236000 358148
rect 236052 358136 236058 358148
rect 399202 358136 399208 358148
rect 236052 358108 399208 358136
rect 236052 358096 236058 358108
rect 399202 358096 399208 358108
rect 399260 358136 399266 358148
rect 399260 358108 402974 358136
rect 399260 358096 399266 358108
rect 38470 358028 38476 358080
rect 38528 358068 38534 358080
rect 200114 358068 200120 358080
rect 38528 358040 200120 358068
rect 38528 358028 38534 358040
rect 200114 358028 200120 358040
rect 200172 358028 200178 358080
rect 216122 358028 216128 358080
rect 216180 358068 216186 358080
rect 227806 358068 227812 358080
rect 216180 358040 227812 358068
rect 216180 358028 216186 358040
rect 227806 358028 227812 358040
rect 227864 358028 227870 358080
rect 396994 358068 397000 358080
rect 238726 358040 397000 358068
rect 216306 357960 216312 358012
rect 216364 358000 216370 358012
rect 231854 358000 231860 358012
rect 216364 357972 231860 358000
rect 216364 357960 216370 357972
rect 231854 357960 231860 357972
rect 231912 357960 231918 358012
rect 218698 357892 218704 357944
rect 218756 357932 218762 357944
rect 230014 357932 230020 357944
rect 218756 357904 230020 357932
rect 218756 357892 218762 357904
rect 230014 357892 230020 357904
rect 230072 357932 230078 357944
rect 238726 357932 238754 358040
rect 396994 358028 397000 358040
rect 397052 358028 397058 358080
rect 402946 358068 402974 358108
rect 416038 358068 416044 358080
rect 402946 358040 416044 358068
rect 416038 358028 416044 358040
rect 416096 358028 416102 358080
rect 308398 357960 308404 358012
rect 308456 358000 308462 358012
rect 359366 358000 359372 358012
rect 308456 357972 359372 358000
rect 308456 357960 308462 357972
rect 359366 357960 359372 357972
rect 359424 357960 359430 358012
rect 230072 357904 238754 357932
rect 230072 357892 230078 357904
rect 311342 357892 311348 357944
rect 311400 357932 311406 357944
rect 356974 357932 356980 357944
rect 311400 357904 356980 357932
rect 311400 357892 311406 357904
rect 356974 357892 356980 357904
rect 357032 357892 357038 357944
rect 218882 357824 218888 357876
rect 218940 357864 218946 357876
rect 223390 357864 223396 357876
rect 218940 357836 223396 357864
rect 218940 357824 218946 357836
rect 223390 357824 223396 357836
rect 223448 357824 223454 357876
rect 314654 357824 314660 357876
rect 314712 357864 314718 357876
rect 358998 357864 359004 357876
rect 314712 357836 359004 357864
rect 314712 357824 314718 357836
rect 358998 357824 359004 357836
rect 359056 357824 359062 357876
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 36538 357456 36544 357468
rect 3384 357428 36544 357456
rect 3384 357416 3390 357428
rect 36538 357416 36544 357428
rect 36596 357416 36602 357468
rect 262122 357348 262128 357400
rect 262180 357388 262186 357400
rect 399294 357388 399300 357400
rect 262180 357360 399300 357388
rect 262180 357348 262186 357360
rect 399294 357348 399300 357360
rect 399352 357388 399358 357400
rect 423122 357388 423128 357400
rect 399352 357360 423128 357388
rect 399352 357348 399358 357360
rect 423122 357348 423128 357360
rect 423180 357388 423186 357400
rect 423582 357388 423588 357400
rect 423180 357360 423588 357388
rect 423180 357348 423186 357360
rect 423582 357348 423588 357360
rect 423640 357348 423646 357400
rect 262766 357280 262772 357332
rect 262824 357320 262830 357332
rect 398190 357320 398196 357332
rect 262824 357292 398196 357320
rect 262824 357280 262830 357292
rect 398190 357280 398196 357292
rect 398248 357320 398254 357332
rect 398650 357320 398656 357332
rect 398248 357292 398656 357320
rect 398248 357280 398254 357292
rect 398650 357280 398656 357292
rect 398708 357280 398714 357332
rect 398834 357280 398840 357332
rect 398892 357320 398898 357332
rect 399110 357320 399116 357332
rect 398892 357292 399116 357320
rect 398892 357280 398898 357292
rect 399110 357280 399116 357292
rect 399168 357320 399174 357332
rect 433426 357320 433432 357332
rect 399168 357292 433432 357320
rect 399168 357280 399174 357292
rect 433426 357280 433432 357292
rect 433484 357320 433490 357332
rect 433484 357292 441614 357320
rect 433484 357280 433490 357292
rect 263594 357212 263600 357264
rect 263652 357252 263658 357264
rect 263962 357252 263968 357264
rect 263652 357224 263968 357252
rect 263652 357212 263658 357224
rect 263962 357212 263968 357224
rect 264020 357252 264026 357264
rect 394234 357252 394240 357264
rect 264020 357224 394240 357252
rect 264020 357212 264026 357224
rect 394234 357212 394240 357224
rect 394292 357212 394298 357264
rect 268286 357144 268292 357196
rect 268344 357184 268350 357196
rect 268562 357184 268568 357196
rect 268344 357156 268568 357184
rect 268344 357144 268350 357156
rect 268562 357144 268568 357156
rect 268620 357184 268626 357196
rect 397362 357184 397368 357196
rect 268620 357156 397368 357184
rect 268620 357144 268626 357156
rect 397362 357144 397368 357156
rect 397420 357144 397426 357196
rect 399018 357144 399024 357196
rect 399076 357184 399082 357196
rect 434622 357184 434628 357196
rect 399076 357156 434628 357184
rect 399076 357144 399082 357156
rect 434622 357144 434628 357156
rect 434680 357144 434686 357196
rect 441586 357184 441614 357292
rect 444282 357212 444288 357264
rect 444340 357252 444346 357264
rect 456794 357252 456800 357264
rect 444340 357224 456800 357252
rect 444340 357212 444346 357224
rect 456794 357212 456800 357224
rect 456852 357212 456858 357264
rect 451458 357184 451464 357196
rect 441586 357156 451464 357184
rect 451458 357144 451464 357156
rect 451516 357144 451522 357196
rect 394050 357076 394056 357128
rect 394108 357116 394114 357128
rect 394418 357116 394424 357128
rect 394108 357088 394424 357116
rect 394108 357076 394114 357088
rect 394418 357076 394424 357088
rect 394476 357116 394482 357128
rect 436002 357116 436008 357128
rect 394476 357088 436008 357116
rect 394476 357076 394482 357088
rect 436002 357076 436008 357088
rect 436060 357076 436066 357128
rect 445662 357076 445668 357128
rect 445720 357116 445726 357128
rect 458174 357116 458180 357128
rect 445720 357088 458180 357116
rect 445720 357076 445726 357088
rect 458174 357076 458180 357088
rect 458232 357076 458238 357128
rect 266354 357008 266360 357060
rect 266412 357048 266418 357060
rect 267550 357048 267556 357060
rect 266412 357020 267556 357048
rect 266412 357008 266418 357020
rect 267550 357008 267556 357020
rect 267608 357048 267614 357060
rect 394602 357048 394608 357060
rect 267608 357020 394608 357048
rect 267608 357008 267614 357020
rect 394602 357008 394608 357020
rect 394660 357048 394666 357060
rect 394660 357020 396396 357048
rect 394660 357008 394666 357020
rect 243538 356940 243544 356992
rect 243596 356980 243602 356992
rect 262122 356980 262128 356992
rect 243596 356952 262128 356980
rect 243596 356940 243602 356952
rect 262122 356940 262128 356952
rect 262180 356940 262186 356992
rect 265066 356940 265072 356992
rect 265124 356980 265130 356992
rect 265710 356980 265716 356992
rect 265124 356952 265716 356980
rect 265124 356940 265130 356952
rect 265710 356940 265716 356952
rect 265768 356980 265774 356992
rect 396368 356980 396396 357020
rect 398374 357008 398380 357060
rect 398432 357048 398438 357060
rect 398742 357048 398748 357060
rect 398432 357020 398748 357048
rect 398432 357008 398438 357020
rect 398742 357008 398748 357020
rect 398800 357048 398806 357060
rect 431954 357048 431960 357060
rect 398800 357020 431960 357048
rect 398800 357008 398806 357020
rect 431954 357008 431960 357020
rect 432012 357048 432018 357060
rect 449986 357048 449992 357060
rect 432012 357020 449992 357048
rect 432012 357008 432018 357020
rect 449986 357008 449992 357020
rect 450044 357008 450050 357060
rect 428550 356980 428556 356992
rect 265768 356952 393314 356980
rect 396368 356952 428556 356980
rect 265768 356940 265774 356952
rect 257338 356872 257344 356924
rect 257396 356912 257402 356924
rect 275922 356912 275928 356924
rect 257396 356884 275928 356912
rect 257396 356872 257402 356884
rect 275922 356872 275928 356884
rect 275980 356872 275986 356924
rect 393286 356912 393314 356952
rect 428550 356940 428556 356952
rect 428608 356940 428614 356992
rect 436002 356940 436008 356992
rect 436060 356980 436066 356992
rect 454034 356980 454040 356992
rect 436060 356952 454040 356980
rect 436060 356940 436066 356952
rect 454034 356940 454040 356952
rect 454092 356940 454098 356992
rect 394326 356912 394332 356924
rect 393286 356884 394332 356912
rect 394326 356872 394332 356884
rect 394384 356912 394390 356924
rect 394602 356912 394608 356924
rect 394384 356884 394608 356912
rect 394384 356872 394390 356884
rect 394602 356872 394608 356884
rect 394660 356872 394666 356924
rect 397270 356872 397276 356924
rect 397328 356912 397334 356924
rect 430666 356912 430672 356924
rect 397328 356884 430672 356912
rect 397328 356872 397334 356884
rect 430666 356872 430672 356884
rect 430724 356872 430730 356924
rect 434622 356872 434628 356924
rect 434680 356912 434686 356924
rect 452746 356912 452752 356924
rect 434680 356884 452752 356912
rect 434680 356872 434686 356884
rect 452746 356872 452752 356884
rect 452804 356872 452810 356924
rect 491938 356872 491944 356924
rect 491996 356912 492002 356924
rect 498194 356912 498200 356924
rect 491996 356884 498200 356912
rect 491996 356872 492002 356884
rect 498194 356872 498200 356884
rect 498252 356872 498258 356924
rect 251266 356804 251272 356856
rect 251324 356844 251330 356856
rect 269758 356844 269764 356856
rect 251324 356816 269764 356844
rect 251324 356804 251330 356816
rect 269758 356804 269764 356816
rect 269816 356844 269822 356856
rect 270402 356844 270408 356856
rect 269816 356816 270408 356844
rect 269816 356804 269822 356816
rect 270402 356804 270408 356816
rect 270460 356804 270466 356856
rect 272150 356804 272156 356856
rect 272208 356844 272214 356856
rect 398834 356844 398840 356856
rect 272208 356816 398840 356844
rect 272208 356804 272214 356816
rect 398834 356804 398840 356816
rect 398892 356804 398898 356856
rect 436830 356804 436836 356856
rect 436888 356844 436894 356856
rect 455414 356844 455420 356856
rect 436888 356816 455420 356844
rect 436888 356804 436894 356816
rect 455414 356804 455420 356816
rect 455472 356804 455478 356856
rect 249702 356736 249708 356788
rect 249760 356776 249766 356788
rect 266354 356776 266360 356788
rect 249760 356748 266360 356776
rect 249760 356736 249766 356748
rect 266354 356736 266360 356748
rect 266412 356736 266418 356788
rect 266446 356736 266452 356788
rect 266504 356776 266510 356788
rect 394510 356776 394516 356788
rect 266504 356748 394516 356776
rect 266504 356736 266510 356748
rect 394510 356736 394516 356748
rect 394568 356776 394574 356788
rect 394568 356748 427308 356776
rect 394568 356736 394574 356748
rect 252094 356668 252100 356720
rect 252152 356708 252158 356720
rect 254578 356708 254584 356720
rect 252152 356680 254584 356708
rect 252152 356668 252158 356680
rect 254578 356668 254584 356680
rect 254636 356708 254642 356720
rect 273346 356708 273352 356720
rect 254636 356680 273352 356708
rect 254636 356668 254642 356680
rect 273346 356668 273352 356680
rect 273404 356708 273410 356720
rect 274450 356708 274456 356720
rect 273404 356680 274456 356708
rect 273404 356668 273410 356680
rect 274450 356668 274456 356680
rect 274508 356668 274514 356720
rect 398190 356668 398196 356720
rect 398248 356708 398254 356720
rect 424962 356708 424968 356720
rect 398248 356680 424968 356708
rect 398248 356668 398254 356680
rect 424962 356668 424968 356680
rect 425020 356668 425026 356720
rect 60642 356600 60648 356652
rect 60700 356640 60706 356652
rect 62758 356640 62764 356652
rect 60700 356612 62764 356640
rect 60700 356600 60706 356612
rect 62758 356600 62764 356612
rect 62816 356600 62822 356652
rect 244918 356600 244924 356652
rect 244976 356640 244982 356652
rect 262766 356640 262772 356652
rect 244976 356612 262772 356640
rect 244976 356600 244982 356612
rect 262766 356600 262772 356612
rect 262824 356600 262830 356652
rect 274542 356600 274548 356652
rect 274600 356640 274606 356652
rect 394418 356640 394424 356652
rect 274600 356612 394424 356640
rect 274600 356600 274606 356612
rect 394418 356600 394424 356612
rect 394476 356600 394482 356652
rect 394602 356600 394608 356652
rect 394660 356640 394666 356652
rect 426894 356640 426900 356652
rect 394660 356612 426900 356640
rect 394660 356600 394666 356612
rect 426894 356600 426900 356612
rect 426952 356600 426958 356652
rect 250070 356532 250076 356584
rect 250128 356572 250134 356584
rect 268286 356572 268292 356584
rect 250128 356544 268292 356572
rect 250128 356532 250134 356544
rect 268286 356532 268292 356544
rect 268344 356532 268350 356584
rect 275922 356532 275928 356584
rect 275980 356572 275986 356584
rect 394142 356572 394148 356584
rect 275980 356544 394148 356572
rect 275980 356532 275986 356544
rect 394142 356532 394148 356544
rect 394200 356532 394206 356584
rect 394234 356532 394240 356584
rect 394292 356572 394298 356584
rect 425422 356572 425428 356584
rect 394292 356544 425428 356572
rect 394292 356532 394298 356544
rect 425422 356532 425428 356544
rect 425480 356572 425486 356584
rect 426342 356572 426348 356584
rect 425480 356544 426348 356572
rect 425480 356532 425486 356544
rect 426342 356532 426348 356544
rect 426400 356532 426406 356584
rect 427280 356572 427308 356748
rect 437566 356736 437572 356788
rect 437624 356776 437630 356788
rect 438394 356776 438400 356788
rect 437624 356748 438400 356776
rect 437624 356736 437630 356748
rect 438394 356736 438400 356748
rect 438452 356776 438458 356788
rect 456794 356776 456800 356788
rect 438452 356748 456800 356776
rect 438452 356736 438458 356748
rect 456794 356736 456800 356748
rect 456852 356736 456858 356788
rect 429194 356668 429200 356720
rect 429252 356708 429258 356720
rect 430022 356708 430028 356720
rect 429252 356680 430028 356708
rect 429252 356668 429258 356680
rect 430022 356668 430028 356680
rect 430080 356708 430086 356720
rect 448514 356708 448520 356720
rect 430080 356680 448520 356708
rect 430080 356668 430086 356680
rect 448514 356668 448520 356680
rect 448572 356668 448578 356720
rect 428550 356600 428556 356652
rect 428608 356640 428614 356652
rect 447134 356640 447140 356652
rect 428608 356612 447140 356640
rect 428608 356600 428614 356612
rect 447134 356600 447140 356612
rect 447192 356600 447198 356652
rect 464430 356600 464436 356652
rect 464488 356640 464494 356652
rect 467834 356640 467840 356652
rect 464488 356612 467840 356640
rect 464488 356600 464494 356612
rect 467834 356600 467840 356612
rect 467892 356600 467898 356652
rect 427630 356572 427636 356584
rect 427280 356544 427636 356572
rect 427630 356532 427636 356544
rect 427688 356572 427694 356584
rect 445754 356572 445760 356584
rect 427688 356544 445760 356572
rect 427688 356532 427694 356544
rect 445754 356532 445760 356544
rect 445812 356532 445818 356584
rect 258810 356464 258816 356516
rect 258868 356504 258874 356516
rect 277026 356504 277032 356516
rect 258868 356476 277032 356504
rect 258868 356464 258874 356476
rect 277026 356464 277032 356476
rect 277084 356504 277090 356516
rect 393774 356504 393780 356516
rect 277084 356476 393780 356504
rect 277084 356464 277090 356476
rect 393774 356464 393780 356476
rect 393832 356504 393838 356516
rect 394602 356504 394608 356516
rect 393832 356476 394608 356504
rect 393832 356464 393838 356476
rect 394602 356464 394608 356476
rect 394660 356464 394666 356516
rect 423582 356464 423588 356516
rect 423640 356504 423646 356516
rect 441706 356504 441712 356516
rect 423640 356476 441712 356504
rect 423640 356464 423646 356476
rect 441706 356464 441712 356476
rect 441764 356464 441770 356516
rect 471238 356464 471244 356516
rect 471296 356504 471302 356516
rect 477494 356504 477500 356516
rect 471296 356476 477500 356504
rect 471296 356464 471302 356476
rect 477494 356464 477500 356476
rect 477552 356464 477558 356516
rect 255314 356396 255320 356448
rect 255372 356436 255378 356448
rect 255774 356436 255780 356448
rect 255372 356408 255780 356436
rect 255372 356396 255378 356408
rect 255774 356396 255780 356408
rect 255832 356436 255838 356448
rect 274542 356436 274548 356448
rect 255832 356408 274548 356436
rect 255832 356396 255838 356408
rect 274542 356396 274548 356408
rect 274600 356396 274606 356448
rect 397362 356396 397368 356448
rect 397420 356436 397426 356448
rect 429194 356436 429200 356448
rect 397420 356408 429200 356436
rect 397420 356396 397426 356408
rect 429194 356396 429200 356408
rect 429252 356396 429258 356448
rect 430666 356396 430672 356448
rect 430724 356436 430730 356448
rect 448514 356436 448520 356448
rect 430724 356408 448520 356436
rect 430724 356396 430730 356408
rect 448514 356396 448520 356408
rect 448572 356396 448578 356448
rect 251450 356328 251456 356380
rect 251508 356368 251514 356380
rect 252278 356368 252284 356380
rect 251508 356340 252284 356368
rect 251508 356328 251514 356340
rect 252278 356328 252284 356340
rect 252336 356368 252342 356380
rect 271138 356368 271144 356380
rect 252336 356340 271144 356368
rect 252336 356328 252342 356340
rect 271138 356328 271144 356340
rect 271196 356368 271202 356380
rect 398374 356368 398380 356380
rect 271196 356340 398380 356368
rect 271196 356328 271202 356340
rect 398374 356328 398380 356340
rect 398432 356328 398438 356380
rect 426342 356328 426348 356380
rect 426400 356368 426406 356380
rect 442994 356368 443000 356380
rect 426400 356340 443000 356368
rect 426400 356328 426406 356340
rect 442994 356328 443000 356340
rect 443052 356328 443058 356380
rect 479518 356328 479524 356380
rect 479576 356368 479582 356380
rect 488534 356368 488540 356380
rect 479576 356340 488540 356368
rect 479576 356328 479582 356340
rect 488534 356328 488540 356340
rect 488592 356328 488598 356380
rect 77202 356260 77208 356312
rect 77260 356300 77266 356312
rect 196526 356300 196532 356312
rect 77260 356272 196532 356300
rect 77260 356260 77266 356272
rect 196526 356260 196532 356272
rect 196584 356260 196590 356312
rect 244274 356260 244280 356312
rect 244332 356300 244338 356312
rect 245562 356300 245568 356312
rect 244332 356272 245568 356300
rect 244332 356260 244338 356272
rect 245562 356260 245568 356272
rect 245620 356300 245626 356312
rect 263594 356300 263600 356312
rect 245620 356272 263600 356300
rect 245620 356260 245626 356272
rect 263594 356260 263600 356272
rect 263652 356260 263658 356312
rect 270402 356260 270408 356312
rect 270460 356300 270466 356312
rect 397270 356300 397276 356312
rect 270460 356272 397276 356300
rect 270460 356260 270466 356272
rect 397270 356260 397276 356272
rect 397328 356260 397334 356312
rect 426894 356260 426900 356312
rect 426952 356300 426958 356312
rect 444374 356300 444380 356312
rect 426952 356272 444380 356300
rect 426952 356260 426958 356272
rect 444374 356260 444380 356272
rect 444432 356260 444438 356312
rect 467190 356260 467196 356312
rect 467248 356300 467254 356312
rect 474734 356300 474740 356312
rect 467248 356272 474740 356300
rect 467248 356260 467254 356272
rect 474734 356260 474740 356272
rect 474792 356260 474798 356312
rect 476758 356260 476764 356312
rect 476816 356300 476822 356312
rect 483014 356300 483020 356312
rect 476816 356272 483020 356300
rect 476816 356260 476822 356272
rect 483014 356260 483020 356272
rect 483072 356260 483078 356312
rect 494698 356260 494704 356312
rect 494756 356300 494762 356312
rect 500954 356300 500960 356312
rect 494756 356272 500960 356300
rect 494756 356260 494762 356272
rect 500954 356260 500960 356272
rect 501012 356260 501018 356312
rect 68922 356192 68928 356244
rect 68980 356232 68986 356244
rect 192110 356232 192116 356244
rect 68980 356204 192116 356232
rect 68980 356192 68986 356204
rect 192110 356192 192116 356204
rect 192168 356192 192174 356244
rect 245654 356192 245660 356244
rect 245712 356232 245718 356244
rect 246850 356232 246856 356244
rect 245712 356204 246856 356232
rect 245712 356192 245718 356204
rect 246850 356192 246856 356204
rect 246908 356232 246914 356244
rect 265066 356232 265072 356244
rect 246908 356204 265072 356232
rect 246908 356192 246914 356204
rect 265066 356192 265072 356204
rect 265124 356192 265130 356244
rect 274450 356192 274456 356244
rect 274508 356232 274514 356244
rect 399018 356232 399024 356244
rect 274508 356204 399024 356232
rect 274508 356192 274514 356204
rect 399018 356192 399024 356204
rect 399076 356192 399082 356244
rect 424962 356192 424968 356244
rect 425020 356232 425026 356244
rect 441982 356232 441988 356244
rect 425020 356204 441988 356232
rect 425020 356192 425026 356204
rect 441982 356192 441988 356204
rect 442040 356192 442046 356244
rect 482278 356192 482284 356244
rect 482336 356232 482342 356244
rect 489914 356232 489920 356244
rect 482336 356204 489920 356232
rect 482336 356192 482342 356204
rect 489914 356192 489920 356204
rect 489972 356192 489978 356244
rect 74074 356124 74080 356176
rect 74132 356164 74138 356176
rect 203150 356164 203156 356176
rect 74132 356136 203156 356164
rect 74132 356124 74138 356136
rect 203150 356124 203156 356136
rect 203208 356124 203214 356176
rect 233694 356124 233700 356176
rect 233752 356164 233758 356176
rect 248690 356164 248696 356176
rect 233752 356136 248696 356164
rect 233752 356124 233758 356136
rect 248690 356124 248696 356136
rect 248748 356164 248754 356176
rect 249702 356164 249708 356176
rect 248748 356136 249708 356164
rect 248748 356124 248754 356136
rect 249702 356124 249708 356136
rect 249760 356124 249766 356176
rect 252830 356124 252836 356176
rect 252888 356164 252894 356176
rect 253382 356164 253388 356176
rect 252888 356136 253388 356164
rect 252888 356124 252894 356136
rect 253382 356124 253388 356136
rect 253440 356164 253446 356176
rect 272150 356164 272156 356176
rect 253440 356136 272156 356164
rect 253440 356124 253446 356136
rect 272150 356124 272156 356136
rect 272208 356124 272214 356176
rect 394142 356124 394148 356176
rect 394200 356164 394206 356176
rect 436830 356164 436836 356176
rect 394200 356136 436836 356164
rect 394200 356124 394206 356136
rect 436830 356124 436836 356136
rect 436888 356124 436894 356176
rect 472710 356124 472716 356176
rect 472768 356164 472774 356176
rect 480530 356164 480536 356176
rect 472768 356136 480536 356164
rect 472768 356124 472774 356136
rect 480530 356124 480536 356136
rect 480588 356124 480594 356176
rect 487798 356124 487804 356176
rect 487856 356164 487862 356176
rect 495434 356164 495440 356176
rect 487856 356136 495440 356164
rect 487856 356124 487862 356136
rect 495434 356124 495440 356136
rect 495492 356124 495498 356176
rect 64322 356056 64328 356108
rect 64380 356096 64386 356108
rect 65518 356096 65524 356108
rect 64380 356068 65524 356096
rect 64380 356056 64386 356068
rect 65518 356056 65524 356068
rect 65576 356056 65582 356108
rect 68922 356056 68928 356108
rect 68980 356096 68986 356108
rect 198366 356096 198372 356108
rect 68980 356068 198372 356096
rect 68980 356056 68986 356068
rect 198366 356056 198372 356068
rect 198424 356056 198430 356108
rect 247126 356056 247132 356108
rect 247184 356096 247190 356108
rect 266446 356096 266452 356108
rect 247184 356068 266452 356096
rect 247184 356056 247190 356068
rect 266446 356056 266452 356068
rect 266504 356056 266510 356108
rect 394602 356056 394608 356108
rect 394660 356096 394666 356108
rect 437566 356096 437572 356108
rect 394660 356068 437572 356096
rect 394660 356056 394666 356068
rect 437566 356056 437572 356068
rect 437624 356056 437630 356108
rect 457438 356056 457444 356108
rect 457496 356096 457502 356108
rect 460934 356096 460940 356108
rect 457496 356068 460940 356096
rect 457496 356056 457502 356068
rect 460934 356056 460940 356068
rect 460992 356056 460998 356108
rect 467098 356056 467104 356108
rect 467156 356096 467162 356108
rect 470778 356096 470784 356108
rect 467156 356068 470784 356096
rect 467156 356056 467162 356068
rect 470778 356056 470784 356068
rect 470836 356056 470842 356108
rect 476850 356056 476856 356108
rect 476908 356096 476914 356108
rect 492674 356096 492680 356108
rect 476908 356068 492680 356096
rect 476908 356056 476914 356068
rect 492674 356056 492680 356068
rect 492732 356056 492738 356108
rect 497458 356056 497464 356108
rect 497516 356096 497522 356108
rect 505094 356096 505100 356108
rect 497516 356068 505100 356096
rect 497516 356056 497522 356068
rect 505094 356056 505100 356068
rect 505152 356056 505158 356108
rect 210510 355988 210516 356040
rect 210568 356028 210574 356040
rect 260190 356028 260196 356040
rect 210568 356000 260196 356028
rect 210568 355988 210574 356000
rect 260190 355988 260196 356000
rect 260248 355988 260254 356040
rect 210694 355920 210700 355972
rect 210752 355960 210758 355972
rect 260098 355960 260104 355972
rect 210752 355932 260104 355960
rect 210752 355920 210758 355932
rect 260098 355920 260104 355932
rect 260156 355920 260162 355972
rect 210602 355852 210608 355904
rect 210660 355892 210666 355904
rect 255314 355892 255320 355904
rect 210660 355864 255320 355892
rect 210660 355852 210666 355864
rect 255314 355852 255320 355864
rect 255372 355852 255378 355904
rect 208302 355784 208308 355836
rect 208360 355824 208366 355836
rect 251450 355824 251456 355836
rect 208360 355796 251456 355824
rect 208360 355784 208366 355796
rect 251450 355784 251456 355796
rect 251508 355784 251514 355836
rect 216398 355716 216404 355768
rect 216456 355756 216462 355768
rect 258810 355756 258816 355768
rect 216456 355728 258816 355756
rect 216456 355716 216462 355728
rect 258810 355716 258816 355728
rect 258868 355716 258874 355768
rect 215110 355648 215116 355700
rect 215168 355688 215174 355700
rect 257338 355688 257344 355700
rect 215168 355660 257344 355688
rect 215168 355648 215174 355660
rect 257338 355648 257344 355660
rect 257396 355648 257402 355700
rect 210786 355580 210792 355632
rect 210844 355620 210850 355632
rect 244274 355620 244280 355632
rect 210844 355592 244280 355620
rect 210844 355580 210850 355592
rect 244274 355580 244280 355592
rect 244332 355580 244338 355632
rect 275646 355580 275652 355632
rect 275704 355620 275710 355632
rect 292574 355620 292580 355632
rect 275704 355592 292580 355620
rect 275704 355580 275710 355592
rect 292574 355580 292580 355592
rect 292632 355580 292638 355632
rect 310974 355580 310980 355632
rect 311032 355620 311038 355632
rect 322934 355620 322940 355632
rect 311032 355592 322940 355620
rect 311032 355580 311038 355592
rect 322934 355580 322940 355592
rect 322992 355580 322998 355632
rect 217594 355512 217600 355564
rect 217652 355552 217658 355564
rect 251266 355552 251272 355564
rect 217652 355524 251272 355552
rect 217652 355512 217658 355524
rect 251266 355512 251272 355524
rect 251324 355512 251330 355564
rect 290734 355512 290740 355564
rect 290792 355552 290798 355564
rect 360194 355552 360200 355564
rect 290792 355524 360200 355552
rect 290792 355512 290798 355524
rect 360194 355512 360200 355524
rect 360252 355512 360258 355564
rect 216490 355444 216496 355496
rect 216548 355484 216554 355496
rect 250070 355484 250076 355496
rect 216548 355456 250076 355484
rect 216548 355444 216554 355456
rect 250070 355444 250076 355456
rect 250128 355444 250134 355496
rect 287790 355444 287796 355496
rect 287848 355484 287854 355496
rect 360286 355484 360292 355496
rect 287848 355456 360292 355484
rect 287848 355444 287854 355456
rect 360286 355444 360292 355456
rect 360344 355444 360350 355496
rect 219250 355376 219256 355428
rect 219308 355416 219314 355428
rect 251082 355416 251088 355428
rect 219308 355388 251088 355416
rect 219308 355376 219314 355388
rect 251082 355376 251088 355388
rect 251140 355376 251146 355428
rect 284846 355376 284852 355428
rect 284904 355416 284910 355428
rect 361666 355416 361672 355428
rect 284904 355388 361672 355416
rect 284904 355376 284910 355388
rect 361666 355376 361672 355388
rect 361724 355376 361730 355428
rect 39022 355308 39028 355360
rect 39080 355348 39086 355360
rect 199838 355348 199844 355360
rect 39080 355320 199844 355348
rect 39080 355308 39086 355320
rect 199838 355308 199844 355320
rect 199896 355308 199902 355360
rect 217778 355308 217784 355360
rect 217836 355348 217842 355360
rect 247126 355348 247132 355360
rect 217836 355320 247132 355348
rect 217836 355308 217842 355320
rect 247126 355308 247132 355320
rect 247184 355308 247190 355360
rect 281902 355308 281908 355360
rect 281960 355348 281966 355360
rect 359274 355348 359280 355360
rect 281960 355320 359280 355348
rect 281960 355308 281966 355320
rect 359274 355308 359280 355320
rect 359332 355308 359338 355360
rect 218790 355240 218796 355292
rect 218848 355280 218854 355292
rect 238110 355280 238116 355292
rect 218848 355252 238116 355280
rect 218848 355240 218854 355252
rect 238110 355240 238116 355252
rect 238168 355240 238174 355292
rect 239582 355240 239588 355292
rect 239640 355280 239646 355292
rect 264974 355280 264980 355292
rect 239640 355252 264980 355280
rect 239640 355240 239646 355252
rect 264974 355240 264980 355252
rect 265032 355240 265038 355292
rect 217410 355172 217416 355224
rect 217468 355212 217474 355224
rect 230382 355212 230388 355224
rect 217468 355184 230388 355212
rect 217468 355172 217474 355184
rect 230382 355172 230388 355184
rect 230440 355172 230446 355224
rect 210418 355104 210424 355156
rect 210476 355144 210482 355156
rect 225230 355144 225236 355156
rect 210476 355116 225236 355144
rect 210476 355104 210482 355116
rect 225230 355104 225236 355116
rect 225288 355104 225294 355156
rect 251082 354696 251088 354748
rect 251140 354736 251146 354748
rect 252830 354736 252836 354748
rect 251140 354708 252836 354736
rect 251140 354696 251146 354708
rect 252830 354696 252836 354708
rect 252888 354696 252894 354748
rect 278958 354628 278964 354680
rect 279016 354668 279022 354680
rect 357986 354668 357992 354680
rect 279016 354640 357992 354668
rect 279016 354628 279022 354640
rect 357986 354628 357992 354640
rect 358044 354628 358050 354680
rect 309502 354560 309508 354612
rect 309560 354600 309566 354612
rect 392946 354600 392952 354612
rect 309560 354572 392952 354600
rect 309560 354560 309566 354572
rect 392946 354560 392952 354572
rect 393004 354560 393010 354612
rect 306558 354492 306564 354544
rect 306616 354532 306622 354544
rect 393038 354532 393044 354544
rect 306616 354504 393044 354532
rect 306616 354492 306622 354504
rect 393038 354492 393044 354504
rect 393096 354492 393102 354544
rect 303614 354424 303620 354476
rect 303672 354464 303678 354476
rect 392394 354464 392400 354476
rect 303672 354436 392400 354464
rect 303672 354424 303678 354436
rect 392394 354424 392400 354436
rect 392452 354424 392458 354476
rect 297726 354356 297732 354408
rect 297784 354396 297790 354408
rect 395890 354396 395896 354408
rect 297784 354368 395896 354396
rect 297784 354356 297790 354368
rect 395890 354356 395896 354368
rect 395948 354356 395954 354408
rect 294782 354288 294788 354340
rect 294840 354328 294846 354340
rect 395982 354328 395988 354340
rect 294840 354300 395988 354328
rect 294840 354288 294846 354300
rect 395982 354288 395988 354300
rect 396040 354288 396046 354340
rect 291838 354220 291844 354272
rect 291896 354260 291902 354272
rect 395798 354260 395804 354272
rect 291896 354232 395804 354260
rect 291896 354220 291902 354232
rect 395798 354220 395804 354232
rect 395856 354220 395862 354272
rect 269758 354152 269764 354204
rect 269816 354192 269822 354204
rect 287054 354192 287060 354204
rect 269816 354164 287060 354192
rect 269816 354152 269822 354164
rect 287054 354152 287060 354164
rect 287112 354152 287118 354204
rect 288894 354152 288900 354204
rect 288952 354192 288958 354204
rect 395706 354192 395712 354204
rect 288952 354164 395712 354192
rect 288952 354152 288958 354164
rect 395706 354152 395712 354164
rect 395764 354152 395770 354204
rect 285950 354084 285956 354136
rect 286008 354124 286014 354136
rect 395614 354124 395620 354136
rect 286008 354096 395620 354124
rect 286008 354084 286014 354096
rect 395614 354084 395620 354096
rect 395672 354084 395678 354136
rect 283006 354016 283012 354068
rect 283064 354056 283070 354068
rect 395430 354056 395436 354068
rect 283064 354028 395436 354056
rect 283064 354016 283070 354028
rect 395430 354016 395436 354028
rect 395488 354016 395494 354068
rect 38838 353948 38844 354000
rect 38896 353988 38902 354000
rect 198734 353988 198740 354000
rect 38896 353960 198740 353988
rect 38896 353948 38902 353960
rect 198734 353948 198740 353960
rect 198792 353948 198798 354000
rect 218422 353948 218428 354000
rect 218480 353988 218486 354000
rect 226334 353988 226340 354000
rect 218480 353960 226340 353988
rect 218480 353948 218486 353960
rect 226334 353948 226340 353960
rect 226392 353948 226398 354000
rect 231486 353948 231492 354000
rect 231544 353988 231550 354000
rect 260834 353988 260840 354000
rect 231544 353960 260840 353988
rect 231544 353948 231550 353960
rect 260834 353948 260840 353960
rect 260892 353948 260898 354000
rect 280062 353948 280068 354000
rect 280120 353988 280126 354000
rect 395522 353988 395528 354000
rect 280120 353960 395528 353988
rect 280120 353948 280126 353960
rect 395522 353948 395528 353960
rect 395580 353948 395586 354000
rect 288158 353880 288164 353932
rect 288216 353920 288222 353932
rect 358906 353920 358912 353932
rect 288216 353892 358912 353920
rect 288216 353880 288222 353892
rect 358906 353880 358912 353892
rect 358964 353880 358970 353932
rect 291102 353812 291108 353864
rect 291160 353852 291166 353864
rect 357434 353852 357440 353864
rect 291160 353824 357440 353852
rect 291160 353812 291166 353824
rect 357434 353812 357440 353824
rect 357492 353812 357498 353864
rect 313918 353744 313924 353796
rect 313976 353784 313982 353796
rect 325694 353784 325700 353796
rect 313976 353756 325700 353784
rect 313976 353744 313982 353756
rect 325694 353744 325700 353756
rect 325752 353744 325758 353796
rect 219802 353200 219808 353252
rect 219860 353240 219866 353252
rect 252094 353240 252100 353252
rect 219860 353212 252100 353240
rect 219860 353200 219866 353212
rect 252094 353200 252100 353212
rect 252152 353200 252158 353252
rect 38930 352520 38936 352572
rect 38988 352560 38994 352572
rect 197630 352560 197636 352572
rect 38988 352532 197636 352560
rect 38988 352520 38994 352532
rect 197630 352520 197636 352532
rect 197688 352520 197694 352572
rect 215754 352520 215760 352572
rect 215812 352560 215818 352572
rect 238754 352560 238760 352572
rect 215812 352532 238760 352560
rect 215812 352520 215818 352532
rect 238754 352520 238760 352532
rect 238812 352520 238818 352572
rect 191190 351908 191196 351960
rect 191248 351948 191254 351960
rect 580166 351948 580172 351960
rect 191248 351920 580172 351948
rect 191248 351908 191254 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 213362 351840 213368 351892
rect 213420 351880 213426 351892
rect 237006 351880 237012 351892
rect 213420 351852 237012 351880
rect 213420 351840 213426 351852
rect 237006 351840 237012 351852
rect 237064 351840 237070 351892
rect 280430 351840 280436 351892
rect 280488 351880 280494 351892
rect 390370 351880 390376 351892
rect 280488 351852 390376 351880
rect 280488 351840 280494 351852
rect 390370 351840 390376 351852
rect 390428 351840 390434 351892
rect 210878 351772 210884 351824
rect 210936 351812 210942 351824
rect 215754 351812 215760 351824
rect 210936 351784 215760 351812
rect 210936 351772 210942 351784
rect 215754 351772 215760 351784
rect 215812 351812 215818 351824
rect 216398 351812 216404 351824
rect 215812 351784 216404 351812
rect 215812 351772 215818 351784
rect 216398 351772 216404 351784
rect 216456 351772 216462 351824
rect 253198 351772 253204 351824
rect 253256 351812 253262 351824
rect 276014 351812 276020 351824
rect 253256 351784 276020 351812
rect 253256 351772 253262 351784
rect 276014 351772 276020 351784
rect 276072 351772 276078 351824
rect 277486 351772 277492 351824
rect 277544 351812 277550 351824
rect 390002 351812 390008 351824
rect 277544 351784 390008 351812
rect 277544 351772 277550 351784
rect 390002 351772 390008 351784
rect 390060 351772 390066 351824
rect 274542 351704 274548 351756
rect 274600 351744 274606 351756
rect 389726 351744 389732 351756
rect 274600 351716 389732 351744
rect 274600 351704 274606 351716
rect 389726 351704 389732 351716
rect 389784 351704 389790 351756
rect 271598 351636 271604 351688
rect 271656 351676 271662 351688
rect 390278 351676 390284 351688
rect 271656 351648 390284 351676
rect 271656 351636 271662 351648
rect 390278 351636 390284 351648
rect 390336 351636 390342 351688
rect 268286 351568 268292 351620
rect 268344 351608 268350 351620
rect 390462 351608 390468 351620
rect 268344 351580 390468 351608
rect 268344 351568 268350 351580
rect 390462 351568 390468 351580
rect 390520 351568 390526 351620
rect 264974 351500 264980 351552
rect 265032 351540 265038 351552
rect 390094 351540 390100 351552
rect 265032 351512 390100 351540
rect 265032 351500 265038 351512
rect 390094 351500 390100 351512
rect 390152 351500 390158 351552
rect 261662 351432 261668 351484
rect 261720 351472 261726 351484
rect 389818 351472 389824 351484
rect 261720 351444 389824 351472
rect 261720 351432 261726 351444
rect 389818 351432 389824 351444
rect 389876 351432 389882 351484
rect 251726 351364 251732 351416
rect 251784 351404 251790 351416
rect 392854 351404 392860 351416
rect 251784 351376 392860 351404
rect 251784 351364 251790 351376
rect 392854 351364 392860 351376
rect 392912 351364 392918 351416
rect 225322 351296 225328 351348
rect 225380 351336 225386 351348
rect 245654 351336 245660 351348
rect 225380 351308 245660 351336
rect 225380 351296 225386 351308
rect 245654 351296 245660 351308
rect 245712 351296 245718 351348
rect 248046 351296 248052 351348
rect 248104 351336 248110 351348
rect 392762 351336 392768 351348
rect 248104 351308 392768 351336
rect 248104 351296 248110 351308
rect 392762 351296 392768 351308
rect 392820 351296 392826 351348
rect 244734 351228 244740 351280
rect 244792 351268 244798 351280
rect 393222 351268 393228 351280
rect 244792 351240 393228 351268
rect 244792 351228 244798 351240
rect 393222 351228 393228 351240
rect 393280 351228 393286 351280
rect 38378 351160 38384 351212
rect 38436 351200 38442 351212
rect 191374 351200 191380 351212
rect 38436 351172 191380 351200
rect 38436 351160 38442 351172
rect 191374 351160 191380 351172
rect 191432 351160 191438 351212
rect 241054 351160 241060 351212
rect 241112 351200 241118 351212
rect 392486 351200 392492 351212
rect 241112 351172 392492 351200
rect 241112 351160 241118 351172
rect 392486 351160 392492 351172
rect 392544 351160 392550 351212
rect 283374 351092 283380 351144
rect 283432 351132 283438 351144
rect 390186 351132 390192 351144
rect 283432 351104 390192 351132
rect 283432 351092 283438 351104
rect 390186 351092 390192 351104
rect 390244 351092 390250 351144
rect 312446 351024 312452 351076
rect 312504 351064 312510 351076
rect 399478 351064 399484 351076
rect 312504 351036 399484 351064
rect 312504 351024 312510 351036
rect 399478 351024 399484 351036
rect 399536 351024 399542 351076
rect 315390 350956 315396 351008
rect 315448 350996 315454 351008
rect 393130 350996 393136 351008
rect 315448 350968 393136 350996
rect 315448 350956 315454 350968
rect 393130 350956 393136 350968
rect 393188 350956 393194 351008
rect 212718 350548 212724 350600
rect 212776 350588 212782 350600
rect 213362 350588 213368 350600
rect 212776 350560 213368 350588
rect 212776 350548 212782 350560
rect 213362 350548 213368 350560
rect 213420 350548 213426 350600
rect 213454 350480 213460 350532
rect 213512 350520 213518 350532
rect 225322 350520 225328 350532
rect 213512 350492 225328 350520
rect 213512 350480 213518 350492
rect 225322 350480 225328 350492
rect 225380 350520 225386 350532
rect 225598 350520 225604 350532
rect 225380 350492 225604 350520
rect 225380 350480 225386 350492
rect 225598 350480 225604 350492
rect 225656 350480 225662 350532
rect 248782 350480 248788 350532
rect 248840 350520 248846 350532
rect 251082 350520 251088 350532
rect 248840 350492 251088 350520
rect 248840 350480 248846 350492
rect 251082 350480 251088 350492
rect 251140 350480 251146 350532
rect 93394 349800 93400 349852
rect 93452 349840 93458 349852
rect 202966 349840 202972 349852
rect 93452 349812 202972 349840
rect 93452 349800 93458 349812
rect 202966 349800 202972 349812
rect 203024 349800 203030 349852
rect 247678 349800 247684 349852
rect 247736 349840 247742 349852
rect 449894 349840 449900 349852
rect 247736 349812 449900 349840
rect 247736 349800 247742 349812
rect 449894 349800 449900 349812
rect 449952 349800 449958 349852
rect 217042 349052 217048 349104
rect 217100 349092 217106 349104
rect 233694 349092 233700 349104
rect 217100 349064 233700 349092
rect 217100 349052 217106 349064
rect 233694 349052 233700 349064
rect 233752 349052 233758 349104
rect 303982 349052 303988 349104
rect 304040 349092 304046 349104
rect 387242 349092 387248 349104
rect 304040 349064 387248 349092
rect 304040 349052 304046 349064
rect 387242 349052 387248 349064
rect 387300 349052 387306 349104
rect 301038 348984 301044 349036
rect 301096 349024 301102 349036
rect 387426 349024 387432 349036
rect 301096 348996 387432 349024
rect 301096 348984 301102 348996
rect 387426 348984 387432 348996
rect 387484 348984 387490 349036
rect 298094 348916 298100 348968
rect 298152 348956 298158 348968
rect 387610 348956 387616 348968
rect 298152 348928 387616 348956
rect 298152 348916 298158 348928
rect 387610 348916 387616 348928
rect 387668 348916 387674 348968
rect 295150 348848 295156 348900
rect 295208 348888 295214 348900
rect 387334 348888 387340 348900
rect 295208 348860 387340 348888
rect 295208 348848 295214 348860
rect 387334 348848 387340 348860
rect 387392 348848 387398 348900
rect 292206 348780 292212 348832
rect 292264 348820 292270 348832
rect 387150 348820 387156 348832
rect 292264 348792 387156 348820
rect 292264 348780 292270 348792
rect 387150 348780 387156 348792
rect 387208 348780 387214 348832
rect 289262 348712 289268 348764
rect 289320 348752 289326 348764
rect 387518 348752 387524 348764
rect 289320 348724 387524 348752
rect 289320 348712 289326 348724
rect 387518 348712 387524 348724
rect 387576 348712 387582 348764
rect 286318 348644 286324 348696
rect 286376 348684 286382 348696
rect 389910 348684 389916 348696
rect 286376 348656 389916 348684
rect 286376 348644 286382 348656
rect 389910 348644 389916 348656
rect 389968 348644 389974 348696
rect 248414 348576 248420 348628
rect 248472 348616 248478 348628
rect 384482 348616 384488 348628
rect 248472 348588 384488 348616
rect 248472 348576 248478 348588
rect 384482 348576 384488 348588
rect 384540 348576 384546 348628
rect 76006 348508 76012 348560
rect 76064 348548 76070 348560
rect 205358 348548 205364 348560
rect 76064 348520 205364 348548
rect 76064 348508 76070 348520
rect 205358 348508 205364 348520
rect 205416 348508 205422 348560
rect 245102 348508 245108 348560
rect 245160 348548 245166 348560
rect 384298 348548 384304 348560
rect 245160 348520 384304 348548
rect 245160 348508 245166 348520
rect 384298 348508 384304 348520
rect 384356 348508 384362 348560
rect 14550 348440 14556 348492
rect 14608 348480 14614 348492
rect 154942 348480 154948 348492
rect 14608 348452 154948 348480
rect 14608 348440 14614 348452
rect 154942 348440 154948 348452
rect 155000 348440 155006 348492
rect 241422 348440 241428 348492
rect 241480 348480 241486 348492
rect 384390 348480 384396 348492
rect 241480 348452 384396 348480
rect 241480 348440 241486 348452
rect 384390 348440 384396 348452
rect 384448 348440 384454 348492
rect 134334 348372 134340 348424
rect 134392 348412 134398 348424
rect 580442 348412 580448 348424
rect 134392 348384 580448 348412
rect 134392 348372 134398 348384
rect 580442 348372 580448 348384
rect 580500 348372 580506 348424
rect 306926 348304 306932 348356
rect 306984 348344 306990 348356
rect 387058 348344 387064 348356
rect 306984 348316 387064 348344
rect 306984 348304 306990 348316
rect 387058 348304 387064 348316
rect 387116 348304 387122 348356
rect 309870 348236 309876 348288
rect 309928 348276 309934 348288
rect 387702 348276 387708 348288
rect 309928 348248 387708 348276
rect 309928 348236 309934 348248
rect 387702 348236 387708 348248
rect 387760 348236 387766 348288
rect 312814 348168 312820 348220
rect 312872 348208 312878 348220
rect 386966 348208 386972 348220
rect 312872 348180 386972 348208
rect 312872 348168 312878 348180
rect 386966 348168 386972 348180
rect 387024 348168 387030 348220
rect 78490 347080 78496 347132
rect 78548 347120 78554 347132
rect 206094 347120 206100 347132
rect 78548 347092 206100 347120
rect 78548 347080 78554 347092
rect 206094 347080 206100 347092
rect 206152 347080 206158 347132
rect 133598 347012 133604 347064
rect 133656 347052 133662 347064
rect 540330 347052 540336 347064
rect 133656 347024 540336 347052
rect 133656 347012 133662 347024
rect 540330 347012 540336 347024
rect 540388 347012 540394 347064
rect 140222 345652 140228 345704
rect 140280 345692 140286 345704
rect 558914 345692 558920 345704
rect 140280 345664 558920 345692
rect 140280 345652 140286 345664
rect 558914 345652 558920 345664
rect 558972 345652 558978 345704
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 148318 345080 148324 345092
rect 3384 345052 148324 345080
rect 3384 345040 3390 345052
rect 148318 345040 148324 345052
rect 148376 345040 148382 345092
rect 212350 344972 212356 345024
rect 212408 345012 212414 345024
rect 243538 345012 243544 345024
rect 212408 344984 243544 345012
rect 212408 344972 212414 344984
rect 243538 344972 243544 344984
rect 243596 344972 243602 345024
rect 211706 344564 211712 344616
rect 211764 344604 211770 344616
rect 212350 344604 212356 344616
rect 211764 344576 212356 344604
rect 211764 344564 211770 344576
rect 212350 344564 212356 344576
rect 212408 344564 212414 344616
rect 73062 344360 73068 344412
rect 73120 344400 73126 344412
rect 202414 344400 202420 344412
rect 73120 344372 202420 344400
rect 73120 344360 73126 344372
rect 202414 344360 202420 344372
rect 202472 344360 202478 344412
rect 244366 344360 244372 344412
rect 244424 344400 244430 344412
rect 447226 344400 447232 344412
rect 244424 344372 447232 344400
rect 244424 344360 244430 344372
rect 447226 344360 447232 344372
rect 447284 344360 447290 344412
rect 136910 344292 136916 344344
rect 136968 344332 136974 344344
rect 537662 344332 537668 344344
rect 136968 344304 537668 344332
rect 136968 344292 136974 344304
rect 537662 344292 537668 344304
rect 537720 344292 537726 344344
rect 257338 342932 257344 342984
rect 257396 342972 257402 342984
rect 258258 342972 258264 342984
rect 257396 342944 258264 342972
rect 257396 342932 257402 342944
rect 258258 342932 258264 342944
rect 258316 342932 258322 342984
rect 38562 342864 38568 342916
rect 38620 342904 38626 342916
rect 207934 342904 207940 342916
rect 38620 342876 207940 342904
rect 38620 342864 38626 342876
rect 207934 342864 207940 342876
rect 207992 342864 207998 342916
rect 228542 342864 228548 342916
rect 228600 342904 228606 342916
rect 437474 342904 437480 342916
rect 228600 342876 437480 342904
rect 228600 342864 228606 342876
rect 437474 342864 437480 342876
rect 437532 342864 437538 342916
rect 213178 342184 213184 342236
rect 213236 342224 213242 342236
rect 238018 342224 238024 342236
rect 213236 342196 238024 342224
rect 213236 342184 213242 342196
rect 238018 342184 238024 342196
rect 238076 342184 238082 342236
rect 81250 341640 81256 341692
rect 81308 341680 81314 341692
rect 207566 341680 207572 341692
rect 81308 341652 207572 341680
rect 81308 341640 81314 341652
rect 207566 341640 207572 341652
rect 207624 341640 207630 341692
rect 237742 341640 237748 341692
rect 237800 341680 237806 341692
rect 250070 341680 250076 341692
rect 237800 341652 250076 341680
rect 237800 341640 237806 341652
rect 250070 341640 250076 341652
rect 250128 341640 250134 341692
rect 18690 341572 18696 341624
rect 18748 341612 18754 341624
rect 150894 341612 150900 341624
rect 18748 341584 150900 341612
rect 18748 341572 18754 341584
rect 150894 341572 150900 341584
rect 150952 341572 150958 341624
rect 236638 341572 236644 341624
rect 236696 341612 236702 341624
rect 443086 341612 443092 341624
rect 236696 341584 443092 341612
rect 236696 341572 236702 341584
rect 443086 341572 443092 341584
rect 443144 341572 443150 341624
rect 142430 341504 142436 341556
rect 142488 341544 142494 341556
rect 392578 341544 392584 341556
rect 142488 341516 392584 341544
rect 142488 341504 142494 341516
rect 392578 341504 392584 341516
rect 392636 341504 392642 341556
rect 211154 340892 211160 340944
rect 211212 340932 211218 340944
rect 213178 340932 213184 340944
rect 211212 340904 213184 340932
rect 211212 340892 211218 340904
rect 213178 340892 213184 340904
rect 213236 340892 213242 340944
rect 216766 340824 216772 340876
rect 216824 340864 216830 340876
rect 217962 340864 217968 340876
rect 216824 340836 217968 340864
rect 216824 340824 216830 340836
rect 217962 340824 217968 340836
rect 218020 340864 218026 340876
rect 244918 340864 244924 340876
rect 218020 340836 244924 340864
rect 218020 340824 218026 340836
rect 244918 340824 244924 340836
rect 244976 340824 244982 340876
rect 36538 340280 36544 340332
rect 36596 340320 36602 340332
rect 157610 340320 157616 340332
rect 36596 340292 157616 340320
rect 36596 340280 36602 340292
rect 157610 340280 157616 340292
rect 157668 340280 157674 340332
rect 77018 340212 77024 340264
rect 77076 340252 77082 340264
rect 204622 340252 204628 340264
rect 77076 340224 204628 340252
rect 77076 340212 77082 340224
rect 204622 340212 204628 340224
rect 204680 340212 204686 340264
rect 227438 340212 227444 340264
rect 227496 340252 227502 340264
rect 258166 340252 258172 340264
rect 227496 340224 258172 340252
rect 227496 340212 227502 340224
rect 258166 340212 258172 340224
rect 258224 340212 258230 340264
rect 139118 340144 139124 340196
rect 139176 340184 139182 340196
rect 538858 340184 538864 340196
rect 139176 340156 538864 340184
rect 139176 340144 139182 340156
rect 538858 340144 538864 340156
rect 538916 340144 538922 340196
rect 139854 338716 139860 338768
rect 139912 338756 139918 338768
rect 580258 338756 580264 338768
rect 139912 338728 580264 338756
rect 139912 338716 139918 338728
rect 580258 338716 580264 338728
rect 580316 338716 580322 338768
rect 224862 337424 224868 337476
rect 224920 337464 224926 337476
rect 395338 337464 395344 337476
rect 224920 337436 395344 337464
rect 224920 337424 224926 337436
rect 395338 337424 395344 337436
rect 395396 337424 395402 337476
rect 61378 337356 61384 337408
rect 61436 337396 61442 337408
rect 195422 337396 195428 337408
rect 61436 337368 195428 337396
rect 61436 337356 61442 337368
rect 195422 337356 195428 337368
rect 195480 337356 195486 337408
rect 250990 337356 250996 337408
rect 251048 337396 251054 337408
rect 452654 337396 452660 337408
rect 251048 337368 452660 337396
rect 251048 337356 251054 337368
rect 452654 337356 452660 337368
rect 452712 337356 452718 337408
rect 7558 335996 7564 336048
rect 7616 336036 7622 336048
rect 154574 336036 154580 336048
rect 7616 336008 154580 336036
rect 7616 335996 7622 336008
rect 154574 335996 154580 336008
rect 154632 335996 154638 336048
rect 240686 335996 240692 336048
rect 240744 336036 240750 336048
rect 445846 336036 445852 336048
rect 240744 336008 445852 336036
rect 240744 335996 240750 336008
rect 445846 335996 445852 336008
rect 445904 335996 445910 336048
rect 4890 333276 4896 333328
rect 4948 333316 4954 333328
rect 152366 333316 152372 333328
rect 4948 333288 152372 333316
rect 4948 333276 4954 333288
rect 152366 333276 152372 333288
rect 152424 333276 152430 333328
rect 141694 333208 141700 333260
rect 141752 333248 141758 333260
rect 360838 333248 360844 333260
rect 141752 333220 360844 333248
rect 141752 333208 141758 333220
rect 360838 333208 360844 333220
rect 360896 333208 360902 333260
rect 4798 331848 4804 331900
rect 4856 331888 4862 331900
rect 151262 331888 151268 331900
rect 4856 331860 151268 331888
rect 4856 331848 4862 331860
rect 151262 331848 151268 331860
rect 151320 331848 151326 331900
rect 224126 331848 224132 331900
rect 224184 331888 224190 331900
rect 434714 331888 434720 331900
rect 224184 331860 434720 331888
rect 224184 331848 224190 331860
rect 434714 331848 434720 331860
rect 434772 331848 434778 331900
rect 63402 330624 63408 330676
rect 63460 330664 63466 330676
rect 192846 330664 192852 330676
rect 63460 330636 192852 330664
rect 63460 330624 63466 330636
rect 192846 330624 192852 330636
rect 192904 330624 192910 330676
rect 223022 330624 223028 330676
rect 223080 330664 223086 330676
rect 255406 330664 255412 330676
rect 223080 330636 255412 330664
rect 223080 330624 223086 330636
rect 255406 330624 255412 330636
rect 255464 330624 255470 330676
rect 3510 330556 3516 330608
rect 3568 330596 3574 330608
rect 156414 330596 156420 330608
rect 3568 330568 156420 330596
rect 3568 330556 3574 330568
rect 156414 330556 156420 330568
rect 156472 330556 156478 330608
rect 215294 330556 215300 330608
rect 215352 330596 215358 330608
rect 430574 330596 430580 330608
rect 215352 330568 430580 330596
rect 215352 330556 215358 330568
rect 430574 330556 430580 330568
rect 430632 330556 430638 330608
rect 143534 330488 143540 330540
rect 143592 330528 143598 330540
rect 364334 330528 364340 330540
rect 143592 330500 364340 330528
rect 143592 330488 143598 330500
rect 364334 330488 364340 330500
rect 364392 330488 364398 330540
rect 70302 329128 70308 329180
rect 70360 329168 70366 329180
rect 200574 329168 200580 329180
rect 70360 329140 200580 329168
rect 70360 329128 70366 329140
rect 200574 329128 200580 329140
rect 200632 329128 200638 329180
rect 284478 329128 284484 329180
rect 284536 329168 284542 329180
rect 300854 329168 300860 329180
rect 284536 329140 300860 329168
rect 284536 329128 284542 329140
rect 300854 329128 300860 329140
rect 300912 329128 300918 329180
rect 14458 329060 14464 329112
rect 14516 329100 14522 329112
rect 153838 329100 153844 329112
rect 14516 329072 153844 329100
rect 14516 329060 14522 329072
rect 153838 329060 153844 329072
rect 153896 329060 153902 329112
rect 210878 329060 210884 329112
rect 210936 329100 210942 329112
rect 427814 329100 427820 329112
rect 210936 329072 427820 329100
rect 210936 329060 210942 329072
rect 427814 329060 427820 329072
rect 427872 329060 427878 329112
rect 68830 327836 68836 327888
rect 68888 327876 68894 327888
rect 199470 327876 199476 327888
rect 68888 327848 199476 327876
rect 68888 327836 68894 327848
rect 199470 327836 199476 327848
rect 199528 327836 199534 327888
rect 214190 327836 214196 327888
rect 214248 327876 214254 327888
rect 249978 327876 249984 327888
rect 214248 327848 249984 327876
rect 214248 327836 214254 327848
rect 249978 327836 249984 327848
rect 250036 327836 250042 327888
rect 11790 327768 11796 327820
rect 11848 327808 11854 327820
rect 156046 327808 156052 327820
rect 11848 327780 156052 327808
rect 11848 327768 11854 327780
rect 156046 327768 156052 327780
rect 156104 327768 156110 327820
rect 232590 327768 232596 327820
rect 232648 327808 232654 327820
rect 440234 327808 440240 327820
rect 232648 327780 440240 327808
rect 232648 327768 232654 327780
rect 440234 327768 440240 327780
rect 440292 327768 440298 327820
rect 133230 327700 133236 327752
rect 133288 327740 133294 327752
rect 542998 327740 543004 327752
rect 133288 327712 543004 327740
rect 133288 327700 133294 327712
rect 542998 327700 543004 327712
rect 543056 327700 543062 327752
rect 59262 326408 59268 326460
rect 59320 326448 59326 326460
rect 192018 326448 192024 326460
rect 59320 326420 192024 326448
rect 59320 326408 59326 326420
rect 192018 326408 192024 326420
rect 192076 326408 192082 326460
rect 138014 326340 138020 326392
rect 138072 326380 138078 326392
rect 538950 326380 538956 326392
rect 138072 326352 538956 326380
rect 138072 326340 138078 326352
rect 538950 326340 538956 326352
rect 539008 326340 539014 326392
rect 143166 324912 143172 324964
rect 143224 324952 143230 324964
rect 366358 324952 366364 324964
rect 143224 324924 366364 324952
rect 143224 324912 143230 324924
rect 366358 324912 366364 324924
rect 366416 324912 366422 324964
rect 131758 324300 131764 324352
rect 131816 324340 131822 324352
rect 580166 324340 580172 324352
rect 131816 324312 580172 324340
rect 131816 324300 131822 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 137646 323688 137652 323740
rect 137704 323728 137710 323740
rect 193858 323728 193864 323740
rect 137704 323700 193864 323728
rect 137704 323688 137710 323700
rect 193858 323688 193864 323700
rect 193916 323688 193922 323740
rect 25590 323620 25596 323672
rect 25648 323660 25654 323672
rect 152734 323660 152740 323672
rect 25648 323632 152740 323660
rect 25648 323620 25654 323632
rect 152734 323620 152740 323632
rect 152792 323620 152798 323672
rect 66162 323552 66168 323604
rect 66220 323592 66226 323604
rect 195790 323592 195796 323604
rect 66220 323564 195796 323592
rect 66220 323552 66226 323564
rect 195790 323552 195796 323564
rect 195848 323552 195854 323604
rect 65518 322260 65524 322312
rect 65576 322300 65582 322312
rect 194318 322300 194324 322312
rect 65576 322272 194324 322300
rect 65576 322260 65582 322272
rect 194318 322260 194324 322272
rect 194376 322260 194382 322312
rect 138382 322192 138388 322244
rect 138440 322232 138446 322244
rect 537478 322232 537484 322244
rect 138440 322204 537484 322232
rect 138440 322192 138446 322204
rect 537478 322192 537484 322204
rect 537536 322192 537542 322244
rect 79962 320900 79968 320952
rect 80020 320940 80026 320952
rect 206830 320940 206836 320952
rect 80020 320912 206836 320940
rect 80020 320900 80026 320912
rect 206830 320900 206836 320912
rect 206888 320900 206894 320952
rect 257614 320900 257620 320952
rect 257672 320940 257678 320952
rect 457530 320940 457536 320952
rect 257672 320912 457536 320940
rect 257672 320900 257678 320912
rect 457530 320900 457536 320912
rect 457588 320900 457594 320952
rect 135070 320832 135076 320884
rect 135128 320872 135134 320884
rect 540238 320872 540244 320884
rect 135128 320844 540244 320872
rect 135128 320832 135134 320844
rect 540238 320832 540244 320844
rect 540296 320832 540302 320884
rect 306190 319472 306196 319524
rect 306248 319512 306254 319524
rect 491938 319512 491944 319524
rect 306248 319484 491944 319512
rect 306248 319472 306254 319484
rect 491938 319472 491944 319484
rect 491996 319472 492002 319524
rect 142062 319404 142068 319456
rect 142120 319444 142126 319456
rect 363598 319444 363604 319456
rect 142120 319416 363604 319444
rect 142120 319404 142126 319416
rect 363598 319404 363604 319416
rect 363656 319404 363662 319456
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 87598 318832 87604 318844
rect 3384 318804 87604 318832
rect 3384 318792 3390 318804
rect 87598 318792 87604 318804
rect 87656 318792 87662 318844
rect 139486 318180 139492 318232
rect 139544 318220 139550 318232
rect 192478 318220 192484 318232
rect 139544 318192 192484 318220
rect 139544 318180 139550 318192
rect 192478 318180 192484 318192
rect 192536 318180 192542 318232
rect 75822 318112 75828 318164
rect 75880 318152 75886 318164
rect 203058 318152 203064 318164
rect 75880 318124 203064 318152
rect 75880 318112 75886 318124
rect 203058 318112 203064 318124
rect 203116 318112 203122 318164
rect 10318 318044 10324 318096
rect 10376 318084 10382 318096
rect 155678 318084 155684 318096
rect 10376 318056 155684 318084
rect 10376 318044 10382 318056
rect 155678 318044 155684 318056
rect 155736 318044 155742 318096
rect 270862 318044 270868 318096
rect 270920 318084 270926 318096
rect 464430 318084 464436 318096
rect 270920 318056 464436 318084
rect 270920 318044 270926 318056
rect 464430 318044 464436 318056
rect 464488 318044 464494 318096
rect 62022 316684 62028 316736
rect 62080 316724 62086 316736
rect 196894 316724 196900 316736
rect 62080 316696 196900 316724
rect 62080 316684 62086 316696
rect 196894 316684 196900 316696
rect 196952 316684 196958 316736
rect 267550 316684 267556 316736
rect 267608 316724 267614 316736
rect 464338 316724 464344 316736
rect 267608 316696 464344 316724
rect 267608 316684 267614 316696
rect 464338 316684 464344 316696
rect 464396 316684 464402 316736
rect 245470 315392 245476 315444
rect 245528 315432 245534 315444
rect 251450 315432 251456 315444
rect 245528 315404 251456 315432
rect 245528 315392 245534 315404
rect 251450 315392 251456 315404
rect 251508 315392 251514 315444
rect 91002 315324 91008 315376
rect 91060 315364 91066 315376
rect 202782 315364 202788 315376
rect 91060 315336 202788 315364
rect 91060 315324 91066 315336
rect 202782 315324 202788 315336
rect 202840 315324 202846 315376
rect 209774 315324 209780 315376
rect 209832 315364 209838 315376
rect 247218 315364 247224 315376
rect 209832 315336 247224 315364
rect 209832 315324 209838 315336
rect 247218 315324 247224 315336
rect 247276 315324 247282 315376
rect 259822 315324 259828 315376
rect 259880 315364 259886 315376
rect 280154 315364 280160 315376
rect 259880 315336 280160 315364
rect 259880 315324 259886 315336
rect 280154 315324 280160 315336
rect 280212 315324 280218 315376
rect 285582 315324 285588 315376
rect 285640 315364 285646 315376
rect 472710 315364 472716 315376
rect 285640 315336 472716 315364
rect 285640 315324 285646 315336
rect 472710 315324 472716 315336
rect 472768 315324 472774 315376
rect 136542 315256 136548 315308
rect 136600 315296 136606 315308
rect 541618 315296 541624 315308
rect 136600 315268 541624 315296
rect 136600 315256 136606 315268
rect 541618 315256 541624 315268
rect 541676 315256 541682 315308
rect 88242 313964 88248 314016
rect 88300 314004 88306 314016
rect 202046 314004 202052 314016
rect 88300 313976 202052 314004
rect 88300 313964 88306 313976
rect 202046 313964 202052 313976
rect 202104 313964 202110 314016
rect 6914 313896 6920 313948
rect 6972 313936 6978 313948
rect 149422 313936 149428 313948
rect 6972 313908 149428 313936
rect 6972 313896 6978 313908
rect 149422 313896 149428 313908
rect 149480 313896 149486 313948
rect 309134 313896 309140 313948
rect 309192 313936 309198 313948
rect 494698 313936 494704 313948
rect 309192 313908 494704 313936
rect 309192 313896 309198 313908
rect 494698 313896 494704 313908
rect 494756 313896 494762 313948
rect 62758 312536 62764 312588
rect 62816 312576 62822 312588
rect 193950 312576 193956 312588
rect 62816 312548 193956 312576
rect 62816 312536 62822 312548
rect 193950 312536 193956 312548
rect 194008 312536 194014 312588
rect 224494 312536 224500 312588
rect 224552 312576 224558 312588
rect 370498 312576 370504 312588
rect 224552 312548 370504 312576
rect 224552 312536 224558 312548
rect 370498 312536 370504 312548
rect 370556 312536 370562 312588
rect 132126 311856 132132 311908
rect 132184 311896 132190 311908
rect 580166 311896 580172 311908
rect 132184 311868 580172 311896
rect 132184 311856 132190 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 78582 311176 78588 311228
rect 78640 311216 78646 311228
rect 197998 311216 198004 311228
rect 78640 311188 198004 311216
rect 78640 311176 78646 311188
rect 197998 311176 198004 311188
rect 198056 311176 198062 311228
rect 31018 311108 31024 311160
rect 31076 311148 31082 311160
rect 150526 311148 150532 311160
rect 31076 311120 150532 311148
rect 31076 311108 31082 311120
rect 150526 311108 150532 311120
rect 150584 311108 150590 311160
rect 300302 311108 300308 311160
rect 300360 311148 300366 311160
rect 476850 311148 476856 311160
rect 300360 311120 476856 311148
rect 300360 311108 300366 311120
rect 476850 311108 476856 311120
rect 476908 311108 476914 311160
rect 81342 309816 81348 309868
rect 81400 309856 81406 309868
rect 199102 309856 199108 309868
rect 81400 309828 199108 309856
rect 81400 309816 81406 309828
rect 199102 309816 199108 309828
rect 199160 309816 199166 309868
rect 15838 309748 15844 309800
rect 15896 309788 15902 309800
rect 155310 309788 155316 309800
rect 15896 309760 155316 309788
rect 15896 309748 15902 309760
rect 155310 309748 155316 309760
rect 155368 309748 155374 309800
rect 303246 309748 303252 309800
rect 303304 309788 303310 309800
rect 487798 309788 487804 309800
rect 303304 309760 487804 309788
rect 303304 309748 303310 309760
rect 487798 309748 487804 309760
rect 487856 309748 487862 309800
rect 35158 308456 35164 308508
rect 35216 308496 35222 308508
rect 153102 308496 153108 308508
rect 35216 308468 153108 308496
rect 35216 308456 35222 308468
rect 153102 308456 153108 308468
rect 153160 308456 153166 308508
rect 74350 308388 74356 308440
rect 74408 308428 74414 308440
rect 195054 308428 195060 308440
rect 74408 308400 195060 308428
rect 74408 308388 74414 308400
rect 195054 308388 195060 308400
rect 195112 308388 195118 308440
rect 279694 308388 279700 308440
rect 279752 308428 279758 308440
rect 467190 308428 467196 308440
rect 279752 308400 467196 308428
rect 279752 308388 279758 308400
rect 467190 308388 467196 308400
rect 467248 308388 467254 308440
rect 106182 307096 106188 307148
rect 106240 307136 106246 307148
rect 207198 307136 207204 307148
rect 106240 307108 207204 307136
rect 106240 307096 106246 307108
rect 207198 307096 207204 307108
rect 207256 307096 207262 307148
rect 8938 307028 8944 307080
rect 8996 307068 9002 307080
rect 153470 307068 153476 307080
rect 8996 307040 153476 307068
rect 8996 307028 9002 307040
rect 153470 307028 153476 307040
rect 153528 307028 153534 307080
rect 243262 307028 243268 307080
rect 243320 307068 243326 307080
rect 267734 307068 267740 307080
rect 243320 307040 267740 307068
rect 243320 307028 243326 307040
rect 267734 307028 267740 307040
rect 267792 307028 267798 307080
rect 282638 307028 282644 307080
rect 282696 307068 282702 307080
rect 471238 307068 471244 307080
rect 282696 307040 471244 307068
rect 282696 307028 282702 307040
rect 471238 307028 471244 307040
rect 471296 307028 471302 307080
rect 137278 305600 137284 305652
rect 137336 305640 137342 305652
rect 188338 305640 188344 305652
rect 137336 305612 188344 305640
rect 137336 305600 137342 305612
rect 188338 305600 188344 305612
rect 188396 305600 188402 305652
rect 254302 305600 254308 305652
rect 254360 305640 254366 305652
rect 454678 305640 454684 305652
rect 254360 305612 454684 305640
rect 254360 305600 254366 305612
rect 454678 305600 454684 305612
rect 454736 305600 454742 305652
rect 3418 304988 3424 305040
rect 3476 305028 3482 305040
rect 90358 305028 90364 305040
rect 3476 305000 90364 305028
rect 3476 304988 3482 305000
rect 90358 304988 90364 305000
rect 90416 304988 90422 305040
rect 256510 304376 256516 304428
rect 256568 304416 256574 304428
rect 277394 304416 277400 304428
rect 256568 304388 277400 304416
rect 256568 304376 256574 304388
rect 277394 304376 277400 304388
rect 277452 304376 277458 304428
rect 235534 304308 235540 304360
rect 235592 304348 235598 304360
rect 263686 304348 263692 304360
rect 235592 304320 263692 304348
rect 235592 304308 235598 304320
rect 263686 304308 263692 304320
rect 263744 304308 263750 304360
rect 278590 304308 278596 304360
rect 278648 304348 278654 304360
rect 295334 304348 295340 304360
rect 278648 304320 295340 304348
rect 278648 304308 278654 304320
rect 295334 304308 295340 304320
rect 295392 304308 295398 304360
rect 104802 304240 104808 304292
rect 104860 304280 104866 304292
rect 206002 304280 206008 304292
rect 104860 304252 206008 304280
rect 104860 304240 104866 304252
rect 206002 304240 206008 304252
rect 206060 304240 206066 304292
rect 260926 304240 260932 304292
rect 260984 304280 260990 304292
rect 457438 304280 457444 304292
rect 260984 304252 457444 304280
rect 260984 304240 260990 304252
rect 457438 304240 457444 304252
rect 457496 304240 457502 304292
rect 102042 302948 102048 303000
rect 102100 302988 102106 303000
rect 205726 302988 205732 303000
rect 102100 302960 205732 302988
rect 102100 302948 102106 302960
rect 205726 302948 205732 302960
rect 205784 302948 205790 303000
rect 11698 302880 11704 302932
rect 11756 302920 11762 302932
rect 151630 302920 151636 302932
rect 11756 302892 151636 302920
rect 11756 302880 11762 302892
rect 151630 302880 151636 302892
rect 151688 302880 151694 302932
rect 288526 302880 288532 302932
rect 288584 302920 288590 302932
rect 476758 302920 476764 302932
rect 288584 302892 476764 302920
rect 288584 302880 288590 302892
rect 476758 302880 476764 302892
rect 476816 302880 476822 302932
rect 99282 301520 99288 301572
rect 99340 301560 99346 301572
rect 204990 301560 204996 301572
rect 99340 301532 204996 301560
rect 99340 301520 99346 301532
rect 204990 301520 204996 301532
rect 205048 301520 205054 301572
rect 26878 301452 26884 301504
rect 26936 301492 26942 301504
rect 149790 301492 149796 301504
rect 26936 301464 149796 301492
rect 26936 301452 26942 301464
rect 149790 301452 149796 301464
rect 149848 301452 149854 301504
rect 276750 301452 276756 301504
rect 276808 301492 276814 301504
rect 472618 301492 472624 301504
rect 276808 301464 472624 301492
rect 276808 301452 276814 301464
rect 472618 301452 472624 301464
rect 472676 301452 472682 301504
rect 96522 300092 96528 300144
rect 96580 300132 96586 300144
rect 204254 300132 204260 300144
rect 96580 300104 204260 300132
rect 96580 300092 96586 300104
rect 204254 300092 204260 300104
rect 204312 300092 204318 300144
rect 273806 300092 273812 300144
rect 273864 300132 273870 300144
rect 467098 300132 467104 300144
rect 273864 300104 467104 300132
rect 273864 300092 273870 300104
rect 467098 300092 467104 300104
rect 467156 300092 467162 300144
rect 258718 299412 258724 299464
rect 258776 299452 258782 299464
rect 262030 299452 262036 299464
rect 258776 299424 262036 299452
rect 258776 299412 258782 299424
rect 262030 299412 262036 299424
rect 262088 299412 262094 299464
rect 71590 298800 71596 298852
rect 71648 298840 71654 298852
rect 193582 298840 193588 298852
rect 71648 298812 193588 298840
rect 71648 298800 71654 298812
rect 193582 298800 193588 298812
rect 193640 298800 193646 298852
rect 25498 298732 25504 298784
rect 25556 298772 25562 298784
rect 151998 298772 152004 298784
rect 25556 298744 152004 298772
rect 25556 298732 25562 298744
rect 151998 298732 152004 298744
rect 152056 298732 152062 298784
rect 258350 298732 258356 298784
rect 258408 298772 258414 298784
rect 356790 298772 356796 298784
rect 258408 298744 356796 298772
rect 258408 298732 258414 298744
rect 356790 298732 356796 298744
rect 356848 298732 356854 298784
rect 131390 298120 131396 298172
rect 131448 298160 131454 298172
rect 580166 298160 580172 298172
rect 131448 298132 580172 298160
rect 131448 298120 131454 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 260190 298052 260196 298104
rect 260248 298092 260254 298104
rect 265342 298092 265348 298104
rect 260248 298064 265348 298092
rect 260248 298052 260254 298064
rect 265342 298052 265348 298064
rect 265400 298052 265406 298104
rect 305086 297712 305092 297764
rect 305144 297752 305150 297764
rect 317414 297752 317420 297764
rect 305144 297724 317420 297752
rect 305144 297712 305150 297724
rect 317414 297712 317420 297724
rect 317472 297712 317478 297764
rect 254670 297644 254676 297696
rect 254728 297684 254734 297696
rect 356698 297684 356704 297696
rect 254728 297656 356704 297684
rect 254728 297644 254734 297656
rect 356698 297644 356704 297656
rect 356756 297644 356762 297696
rect 232958 297576 232964 297628
rect 233016 297616 233022 297628
rect 357066 297616 357072 297628
rect 233016 297588 357072 297616
rect 233016 297576 233022 297588
rect 357066 297576 357072 297588
rect 357124 297576 357130 297628
rect 228910 297508 228916 297560
rect 228968 297548 228974 297560
rect 356882 297548 356888 297560
rect 228968 297520 356888 297548
rect 228968 297508 228974 297520
rect 356882 297508 356888 297520
rect 356940 297508 356946 297560
rect 263134 297440 263140 297492
rect 263192 297480 263198 297492
rect 282914 297480 282920 297492
rect 263192 297452 282920 297480
rect 263192 297440 263198 297452
rect 282914 297440 282920 297452
rect 282972 297440 282978 297492
rect 294414 297440 294420 297492
rect 294472 297480 294478 297492
rect 479518 297480 479524 297492
rect 294472 297452 479524 297480
rect 294472 297440 294478 297452
rect 479518 297440 479524 297452
rect 479576 297440 479582 297492
rect 38746 297372 38752 297424
rect 38804 297412 38810 297424
rect 196158 297412 196164 297424
rect 38804 297384 196164 297412
rect 38804 297372 38810 297384
rect 196158 297372 196164 297384
rect 196216 297372 196222 297424
rect 219710 297372 219716 297424
rect 219768 297412 219774 297424
rect 433334 297412 433340 297424
rect 219768 297384 433340 297412
rect 219768 297372 219774 297384
rect 433334 297372 433340 297384
rect 433392 297372 433398 297424
rect 177942 296216 177948 296268
rect 178000 296256 178006 296268
rect 289998 296256 290004 296268
rect 178000 296228 290004 296256
rect 178000 296216 178006 296228
rect 289998 296216 290004 296228
rect 290056 296216 290062 296268
rect 178954 296148 178960 296200
rect 179012 296188 179018 296200
rect 304718 296188 304724 296200
rect 179012 296160 304724 296188
rect 179012 296148 179018 296160
rect 304718 296148 304724 296160
rect 304776 296148 304782 296200
rect 71682 296080 71688 296132
rect 71740 296120 71746 296132
rect 201862 296120 201868 296132
rect 71740 296092 201868 296120
rect 71740 296080 71746 296092
rect 201862 296080 201868 296092
rect 201920 296080 201926 296132
rect 281534 296080 281540 296132
rect 281592 296120 281598 296132
rect 298186 296120 298192 296132
rect 281592 296092 298192 296120
rect 281592 296080 281598 296092
rect 298186 296080 298192 296092
rect 298244 296080 298250 296132
rect 299198 296080 299204 296132
rect 299256 296120 299262 296132
rect 313274 296120 313280 296132
rect 299256 296092 313280 296120
rect 299256 296080 299262 296092
rect 313274 296080 313280 296092
rect 313332 296080 313338 296132
rect 177206 296012 177212 296064
rect 177264 296052 177270 296064
rect 310606 296052 310612 296064
rect 177264 296024 310612 296052
rect 177264 296012 177270 296024
rect 310606 296012 310612 296024
rect 310664 296012 310670 296064
rect 38654 295944 38660 295996
rect 38712 295984 38718 295996
rect 194686 295984 194692 295996
rect 38712 295956 194692 295984
rect 38712 295944 38718 295956
rect 194686 295944 194692 295956
rect 194744 295944 194750 295996
rect 249886 295944 249892 295996
rect 249944 295984 249950 295996
rect 273346 295984 273352 295996
rect 249944 295956 273352 295984
rect 249944 295944 249950 295956
rect 273346 295944 273352 295956
rect 273404 295944 273410 295996
rect 297358 295944 297364 295996
rect 297416 295984 297422 295996
rect 482278 295984 482284 295996
rect 297416 295956 482284 295984
rect 297416 295944 297422 295956
rect 482278 295944 482284 295956
rect 482336 295944 482342 295996
rect 177850 295060 177856 295112
rect 177908 295100 177914 295112
rect 272334 295100 272340 295112
rect 177908 295072 272340 295100
rect 177908 295060 177914 295072
rect 272334 295060 272340 295072
rect 272392 295060 272398 295112
rect 191098 294992 191104 295044
rect 191156 295032 191162 295044
rect 287054 295032 287060 295044
rect 191156 295004 287060 295032
rect 191156 294992 191162 295004
rect 287054 294992 287060 295004
rect 287112 294992 287118 295044
rect 178678 294924 178684 294976
rect 178736 294964 178742 294976
rect 275278 294964 275284 294976
rect 178736 294936 275284 294964
rect 178736 294924 178742 294936
rect 275278 294924 275284 294936
rect 275336 294924 275342 294976
rect 178862 294856 178868 294908
rect 178920 294896 178926 294908
rect 278222 294896 278228 294908
rect 178920 294868 278228 294896
rect 178920 294856 178926 294868
rect 278222 294856 278228 294868
rect 278280 294856 278286 294908
rect 182818 294788 182824 294840
rect 182876 294828 182882 294840
rect 284110 294828 284116 294840
rect 182876 294800 284116 294828
rect 182876 294788 182882 294800
rect 284110 294788 284116 294800
rect 284168 294788 284174 294840
rect 178770 294720 178776 294772
rect 178828 294760 178834 294772
rect 281166 294760 281172 294772
rect 178828 294732 281172 294760
rect 178828 294720 178834 294732
rect 281166 294720 281172 294732
rect 281224 294720 281230 294772
rect 67542 294652 67548 294704
rect 67600 294692 67606 294704
rect 197262 294692 197268 294704
rect 67600 294664 197268 294692
rect 67600 294652 67606 294664
rect 197262 294652 197268 294664
rect 197320 294652 197326 294704
rect 58618 294584 58624 294636
rect 58676 294624 58682 294636
rect 193214 294624 193220 294636
rect 58676 294596 193220 294624
rect 58676 294584 58682 294596
rect 193214 294584 193220 294596
rect 193272 294584 193278 294636
rect 296254 294584 296260 294636
rect 296312 294624 296318 294636
rect 310514 294624 310520 294636
rect 296312 294596 310520 294624
rect 296312 294584 296318 294596
rect 310514 294584 310520 294596
rect 310572 294584 310578 294636
rect 315022 294584 315028 294636
rect 315080 294624 315086 294636
rect 497458 294624 497464 294636
rect 315080 294596 497464 294624
rect 315080 294584 315086 294596
rect 497458 294584 497464 294596
rect 497516 294584 497522 294636
rect 203978 293904 203984 293956
rect 204036 293944 204042 293956
rect 231118 293944 231124 293956
rect 204036 293916 231124 293944
rect 204036 293904 204042 293916
rect 231118 293904 231124 293916
rect 231176 293904 231182 293956
rect 201034 293836 201040 293888
rect 201092 293876 201098 293888
rect 235166 293876 235172 293888
rect 201092 293848 235172 293876
rect 201092 293836 201098 293848
rect 235166 293836 235172 293848
rect 235224 293836 235230 293888
rect 218606 293768 218612 293820
rect 218664 293808 218670 293820
rect 252646 293808 252652 293820
rect 218664 293780 252652 293808
rect 218664 293768 218670 293780
rect 252646 293768 252652 293780
rect 252704 293768 252710 293820
rect 200850 293700 200856 293752
rect 200908 293740 200914 293752
rect 239214 293740 239220 293752
rect 200908 293712 239220 293740
rect 200908 293700 200914 293712
rect 239214 293700 239220 293712
rect 239272 293700 239278 293752
rect 200942 293632 200948 293684
rect 201000 293672 201006 293684
rect 242894 293672 242900 293684
rect 201000 293644 242900 293672
rect 201000 293632 201006 293644
rect 242894 293632 242900 293644
rect 242952 293632 242958 293684
rect 177758 293564 177764 293616
rect 177816 293604 177822 293616
rect 266078 293604 266084 293616
rect 177816 293576 266084 293604
rect 177816 293564 177822 293576
rect 266078 293564 266084 293576
rect 266136 293564 266142 293616
rect 272702 293564 272708 293616
rect 272760 293604 272766 293616
rect 289906 293604 289912 293616
rect 272760 293576 289912 293604
rect 272760 293564 272766 293576
rect 289906 293564 289912 293576
rect 289964 293564 289970 293616
rect 290366 293564 290372 293616
rect 290424 293604 290430 293616
rect 304994 293604 305000 293616
rect 290424 293576 305000 293604
rect 290424 293564 290430 293576
rect 304994 293564 305000 293576
rect 305052 293564 305058 293616
rect 203702 293496 203708 293548
rect 203760 293536 203766 293548
rect 295886 293536 295892 293548
rect 203760 293508 295892 293536
rect 203760 293496 203766 293508
rect 295886 293496 295892 293508
rect 295944 293496 295950 293548
rect 203794 293428 203800 293480
rect 203852 293468 203858 293480
rect 298830 293468 298836 293480
rect 203852 293440 298836 293468
rect 203852 293428 203858 293440
rect 298830 293428 298836 293440
rect 298888 293428 298894 293480
rect 203886 293360 203892 293412
rect 203944 293400 203950 293412
rect 301774 293400 301780 293412
rect 203944 293372 301780 293400
rect 203944 293360 203950 293372
rect 301774 293360 301780 293372
rect 301832 293360 301838 293412
rect 86862 293292 86868 293344
rect 86920 293332 86926 293344
rect 201310 293332 201316 293344
rect 86920 293304 201316 293332
rect 86920 293292 86926 293304
rect 201310 293292 201316 293304
rect 201368 293292 201374 293344
rect 204070 293292 204076 293344
rect 204128 293332 204134 293344
rect 307662 293332 307668 293344
rect 204128 293304 307668 293332
rect 204128 293292 204134 293304
rect 307662 293292 307668 293304
rect 307720 293292 307726 293344
rect 308030 293292 308036 293344
rect 308088 293332 308094 293344
rect 320174 293332 320180 293344
rect 308088 293304 320180 293332
rect 308088 293292 308094 293304
rect 320174 293292 320180 293304
rect 320232 293292 320238 293344
rect 200758 293224 200764 293276
rect 200816 293264 200822 293276
rect 246206 293264 246212 293276
rect 200816 293236 246212 293264
rect 200816 293224 200822 293236
rect 246206 293224 246212 293236
rect 246264 293224 246270 293276
rect 264238 293224 264244 293276
rect 264296 293264 264302 293276
rect 462314 293264 462320 293276
rect 264296 293236 462320 293264
rect 264296 293224 264302 293236
rect 462314 293224 462320 293236
rect 462372 293224 462378 293276
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 89714 292584 89720 292596
rect 3476 292556 89720 292584
rect 3476 292544 3482 292556
rect 89714 292544 89720 292556
rect 89772 292544 89778 292596
rect 135438 292068 135444 292120
rect 135496 292108 135502 292120
rect 182910 292108 182916 292120
rect 135496 292080 182916 292108
rect 135496 292068 135502 292080
rect 182910 292068 182916 292080
rect 182968 292068 182974 292120
rect 302142 292068 302148 292120
rect 302200 292108 302206 292120
rect 314746 292108 314752 292120
rect 302200 292080 314752 292108
rect 302200 292068 302206 292080
rect 314746 292068 314752 292080
rect 314804 292068 314810 292120
rect 177574 292000 177580 292052
rect 177632 292040 177638 292052
rect 259454 292040 259460 292052
rect 177632 292012 259460 292040
rect 177632 292000 177638 292012
rect 259454 292000 259460 292012
rect 259512 292000 259518 292052
rect 266446 292000 266452 292052
rect 266504 292040 266510 292052
rect 285674 292040 285680 292052
rect 266504 292012 285680 292040
rect 266504 292000 266510 292012
rect 285674 292000 285680 292012
rect 285732 292000 285738 292052
rect 293310 292000 293316 292052
rect 293368 292040 293374 292052
rect 307754 292040 307760 292052
rect 293368 292012 307760 292040
rect 293368 292000 293374 292012
rect 307754 292000 307760 292012
rect 307812 292000 307818 292052
rect 180058 291932 180064 291984
rect 180116 291972 180122 291984
rect 269390 291972 269396 291984
rect 180116 291944 269396 291972
rect 180116 291932 180122 291944
rect 269390 291932 269396 291944
rect 269448 291932 269454 291984
rect 287422 291932 287428 291984
rect 287480 291972 287486 291984
rect 302234 291972 302240 291984
rect 287480 291944 302240 291972
rect 287480 291932 287486 291944
rect 302234 291932 302240 291944
rect 302292 291932 302298 291984
rect 84102 291864 84108 291916
rect 84160 291904 84166 291916
rect 200206 291904 200212 291916
rect 84160 291876 200212 291904
rect 84160 291864 84166 291876
rect 200206 291864 200212 291876
rect 200264 291864 200270 291916
rect 217502 291864 217508 291916
rect 217560 291904 217566 291916
rect 358262 291904 358268 291916
rect 217560 291876 358268 291904
rect 217560 291864 217566 291876
rect 358262 291864 358268 291876
rect 358320 291864 358326 291916
rect 56502 291796 56508 291848
rect 56560 291836 56566 291848
rect 191742 291836 191748 291848
rect 56560 291808 191748 291836
rect 56560 291796 56566 291808
rect 191742 291796 191748 291808
rect 191800 291796 191806 291848
rect 208302 291796 208308 291848
rect 208360 291836 208366 291848
rect 236086 291836 236092 291848
rect 208360 291808 236092 291836
rect 208360 291796 208366 291808
rect 236086 291796 236092 291808
rect 236144 291796 236150 291848
rect 246574 291796 246580 291848
rect 246632 291836 246638 291848
rect 270586 291836 270592 291848
rect 246632 291808 270592 291836
rect 246632 291796 246638 291808
rect 270586 291796 270592 291808
rect 270644 291796 270650 291848
rect 291470 291796 291476 291848
rect 291528 291836 291534 291848
rect 485774 291836 485780 291848
rect 291528 291808 485780 291836
rect 291528 291796 291534 291808
rect 485774 291796 485780 291808
rect 485832 291796 485838 291848
rect 212166 291116 212172 291168
rect 212224 291156 212230 291168
rect 283742 291156 283748 291168
rect 212224 291128 283748 291156
rect 212224 291116 212230 291128
rect 283742 291116 283748 291128
rect 283800 291116 283806 291168
rect 212258 291048 212264 291100
rect 212316 291088 212322 291100
rect 286686 291088 286692 291100
rect 212316 291060 286692 291088
rect 212316 291048 212322 291060
rect 286686 291048 286692 291060
rect 286744 291048 286750 291100
rect 212074 290980 212080 291032
rect 212132 291020 212138 291032
rect 289630 291020 289636 291032
rect 212132 290992 289636 291020
rect 212132 290980 212138 290992
rect 289630 290980 289636 290992
rect 289688 290980 289694 291032
rect 209682 290912 209688 290964
rect 209740 290952 209746 290964
rect 292574 290952 292580 290964
rect 209740 290924 292580 290952
rect 209740 290912 209746 290924
rect 292574 290912 292580 290924
rect 292632 290912 292638 290964
rect 209498 290844 209504 290896
rect 209556 290884 209562 290896
rect 295518 290884 295524 290896
rect 209556 290856 295524 290884
rect 209556 290844 209562 290856
rect 295518 290844 295524 290856
rect 295576 290844 295582 290896
rect 209590 290776 209596 290828
rect 209648 290816 209654 290828
rect 298462 290816 298468 290828
rect 209648 290788 298468 290816
rect 209648 290776 209654 290788
rect 298462 290776 298468 290788
rect 298520 290776 298526 290828
rect 209038 290708 209044 290760
rect 209096 290748 209102 290760
rect 301406 290748 301412 290760
rect 209096 290720 301412 290748
rect 209096 290708 209102 290720
rect 301406 290708 301412 290720
rect 301464 290708 301470 290760
rect 209406 290640 209412 290692
rect 209464 290680 209470 290692
rect 304350 290680 304356 290692
rect 209464 290652 304356 290680
rect 209464 290640 209470 290652
rect 304350 290640 304356 290652
rect 304408 290640 304414 290692
rect 209222 290572 209228 290624
rect 209280 290612 209286 290624
rect 307294 290612 307300 290624
rect 209280 290584 307300 290612
rect 209280 290572 209286 290584
rect 307294 290572 307300 290584
rect 307352 290572 307358 290624
rect 209314 290504 209320 290556
rect 209372 290544 209378 290556
rect 310238 290544 310244 290556
rect 209372 290516 310244 290544
rect 209372 290504 209378 290516
rect 310238 290504 310244 290516
rect 310296 290504 310302 290556
rect 89714 290436 89720 290488
rect 89772 290476 89778 290488
rect 158254 290476 158260 290488
rect 89772 290448 158260 290476
rect 89772 290436 89778 290448
rect 158254 290436 158260 290448
rect 158312 290436 158318 290488
rect 312078 290436 312084 290488
rect 312136 290476 312142 290488
rect 502334 290476 502340 290488
rect 312136 290448 502340 290476
rect 312136 290436 312142 290448
rect 502334 290436 502340 290448
rect 502392 290436 502398 290488
rect 206554 290368 206560 290420
rect 206612 290408 206618 290420
rect 245838 290408 245844 290420
rect 206612 290380 245844 290408
rect 206612 290368 206618 290380
rect 245838 290368 245844 290380
rect 245896 290368 245902 290420
rect 206646 290300 206652 290352
rect 206704 290340 206710 290352
rect 242526 290340 242532 290352
rect 206704 290312 242532 290340
rect 206704 290300 206710 290312
rect 242526 290300 242532 290312
rect 242584 290300 242590 290352
rect 206738 290232 206744 290284
rect 206796 290272 206802 290284
rect 238846 290272 238852 290284
rect 206796 290244 238852 290272
rect 206796 290232 206802 290244
rect 238846 290232 238852 290244
rect 238904 290232 238910 290284
rect 209130 290164 209136 290216
rect 209188 290204 209194 290216
rect 313182 290204 313188 290216
rect 209188 290176 313188 290204
rect 209188 290164 209194 290176
rect 313182 290164 313188 290176
rect 313240 290164 313246 290216
rect 316678 289756 316684 289808
rect 316736 289796 316742 289808
rect 396718 289796 396724 289808
rect 316736 289768 396724 289796
rect 316736 289756 316742 289768
rect 396718 289756 396724 289768
rect 396776 289756 396782 289808
rect 90358 289212 90364 289264
rect 90416 289252 90422 289264
rect 158622 289252 158628 289264
rect 90416 289224 158628 289252
rect 90416 289212 90422 289224
rect 158622 289212 158628 289224
rect 158680 289212 158686 289264
rect 217318 289212 217324 289264
rect 217376 289252 217382 289264
rect 225966 289252 225972 289264
rect 217376 289224 225972 289252
rect 217376 289212 217382 289224
rect 225966 289212 225972 289224
rect 226024 289212 226030 289264
rect 3510 289144 3516 289196
rect 3568 289184 3574 289196
rect 154206 289184 154212 289196
rect 3568 289156 154212 289184
rect 3568 289144 3574 289156
rect 154206 289144 154212 289156
rect 154264 289144 154270 289196
rect 217686 289144 217692 289196
rect 217744 289184 217750 289196
rect 242158 289184 242164 289196
rect 217744 289156 242164 289184
rect 217744 289144 217750 289156
rect 242158 289144 242164 289156
rect 242216 289144 242222 289196
rect 132862 289076 132868 289128
rect 132920 289116 132926 289128
rect 547138 289116 547144 289128
rect 132920 289088 547144 289116
rect 132920 289076 132926 289088
rect 547138 289076 547144 289088
rect 547196 289076 547202 289128
rect 316126 289008 316132 289060
rect 316184 289048 316190 289060
rect 316678 289048 316684 289060
rect 316184 289020 316684 289048
rect 316184 289008 316190 289020
rect 316678 289008 316684 289020
rect 316736 289008 316742 289060
rect 217870 288396 217876 288448
rect 217928 288436 217934 288448
rect 221550 288436 221556 288448
rect 217928 288408 221556 288436
rect 217928 288396 217934 288408
rect 221550 288396 221556 288408
rect 221608 288396 221614 288448
rect 220814 287920 220820 287972
rect 220872 287960 220878 287972
rect 240226 287960 240232 287972
rect 220872 287932 240232 287960
rect 220872 287920 220878 287932
rect 240226 287920 240232 287932
rect 240284 287920 240290 287972
rect 148318 287852 148324 287904
rect 148376 287892 148382 287904
rect 157150 287892 157156 287904
rect 148376 287864 157156 287892
rect 148376 287852 148382 287864
rect 157150 287852 157156 287864
rect 157208 287852 157214 287904
rect 206462 287852 206468 287904
rect 206520 287892 206526 287904
rect 234798 287892 234804 287904
rect 206520 287864 234804 287892
rect 206520 287852 206526 287864
rect 234798 287852 234804 287864
rect 234856 287852 234862 287904
rect 241790 287852 241796 287904
rect 241848 287892 241854 287904
rect 251266 287892 251272 287904
rect 241848 287864 251272 287892
rect 241848 287852 241854 287864
rect 251266 287852 251272 287864
rect 251324 287852 251330 287904
rect 132586 287784 132592 287836
rect 132644 287824 132650 287836
rect 191190 287824 191196 287836
rect 132644 287796 191196 287824
rect 132644 287784 132650 287796
rect 191190 287784 191196 287796
rect 191248 287784 191254 287836
rect 211890 287784 211896 287836
rect 211948 287824 211954 287836
rect 274910 287824 274916 287836
rect 211948 287796 274916 287824
rect 211948 287784 211954 287796
rect 274910 287784 274916 287796
rect 274968 287784 274974 287836
rect 87598 287716 87604 287768
rect 87656 287756 87662 287768
rect 157886 287756 157892 287768
rect 87656 287728 157892 287756
rect 87656 287716 87662 287728
rect 157886 287716 157892 287728
rect 157944 287716 157950 287768
rect 211798 287716 211804 287768
rect 211856 287756 211862 287768
rect 277854 287756 277860 287768
rect 211856 287728 277860 287756
rect 211856 287716 211862 287728
rect 277854 287716 277860 287728
rect 277912 287716 277918 287768
rect 10410 287648 10416 287700
rect 10468 287688 10474 287700
rect 156782 287688 156788 287700
rect 10468 287660 156788 287688
rect 10468 287648 10474 287660
rect 156782 287648 156788 287660
rect 156840 287648 156846 287700
rect 211982 287648 211988 287700
rect 212040 287688 212046 287700
rect 280798 287688 280804 287700
rect 212040 287660 280804 287688
rect 212040 287648 212046 287660
rect 280798 287648 280804 287660
rect 280856 287648 280862 287700
rect 176746 287580 176752 287632
rect 176804 287620 176810 287632
rect 319530 287620 319536 287632
rect 176804 287592 319536 287620
rect 176804 287580 176810 287592
rect 319530 287580 319536 287592
rect 319588 287580 319594 287632
rect 172974 287512 172980 287564
rect 173032 287552 173038 287564
rect 319714 287552 319720 287564
rect 173032 287524 319720 287552
rect 173032 287512 173038 287524
rect 319714 287512 319720 287524
rect 319772 287512 319778 287564
rect 167086 287444 167092 287496
rect 167144 287484 167150 287496
rect 449894 287484 449900 287496
rect 167144 287456 449900 287484
rect 167144 287444 167150 287456
rect 449894 287444 449900 287456
rect 449952 287444 449958 287496
rect 172606 287376 172612 287428
rect 172664 287416 172670 287428
rect 458174 287416 458180 287428
rect 172664 287388 458180 287416
rect 172664 287376 172670 287388
rect 458174 287376 458180 287388
rect 458232 287376 458238 287428
rect 182910 287308 182916 287360
rect 182968 287348 182974 287360
rect 471974 287348 471980 287360
rect 182968 287320 471980 287348
rect 182968 287308 182974 287320
rect 471974 287308 471980 287320
rect 472032 287308 472038 287360
rect 184382 287240 184388 287292
rect 184440 287280 184446 287292
rect 474734 287280 474740 287292
rect 184440 287252 474740 287280
rect 184440 287240 184446 287252
rect 474734 287240 474740 287252
rect 474792 287240 474798 287292
rect 187326 287172 187332 287224
rect 187384 287212 187390 287224
rect 478874 287212 478880 287224
rect 187384 287184 478880 287212
rect 187384 287172 187390 287184
rect 478874 287172 478880 287184
rect 478932 287172 478938 287224
rect 189534 287104 189540 287156
rect 189592 287144 189598 287156
rect 484394 287144 484400 287156
rect 189592 287116 484400 287144
rect 189592 287104 189598 287116
rect 484394 287104 484400 287116
rect 484452 287104 484458 287156
rect 190638 287036 190644 287088
rect 190696 287076 190702 287088
rect 485774 287076 485780 287088
rect 190696 287048 485780 287076
rect 190696 287036 190702 287048
rect 485774 287036 485780 287048
rect 485832 287036 485838 287088
rect 146110 286492 146116 286544
rect 146168 286532 146174 286544
rect 201494 286532 201500 286544
rect 146168 286504 201500 286532
rect 146168 286492 146174 286504
rect 201494 286492 201500 286504
rect 201552 286492 201558 286544
rect 221458 286492 221464 286544
rect 221516 286532 221522 286544
rect 244274 286532 244280 286544
rect 221516 286504 244280 286532
rect 221516 286492 221522 286504
rect 244274 286492 244280 286504
rect 244332 286492 244338 286544
rect 166902 286424 166908 286476
rect 166960 286464 166966 286476
rect 364334 286464 364340 286476
rect 166960 286436 364340 286464
rect 166960 286424 166966 286436
rect 364334 286424 364340 286436
rect 364392 286424 364398 286476
rect 168834 286356 168840 286408
rect 168892 286396 168898 286408
rect 368474 286396 368480 286408
rect 168892 286368 368480 286396
rect 168892 286356 168898 286368
rect 368474 286356 368480 286368
rect 368532 286356 368538 286408
rect 170674 286288 170680 286340
rect 170732 286328 170738 286340
rect 373994 286328 374000 286340
rect 170732 286300 374000 286328
rect 170732 286288 170738 286300
rect 373994 286288 374000 286300
rect 374052 286288 374058 286340
rect 172422 286220 172428 286272
rect 172480 286260 172486 286272
rect 378134 286260 378140 286272
rect 172480 286232 378140 286260
rect 172480 286220 172486 286232
rect 378134 286220 378140 286232
rect 378192 286220 378198 286272
rect 174354 286152 174360 286204
rect 174412 286192 174418 286204
rect 383654 286192 383660 286204
rect 174412 286164 383660 286192
rect 174412 286152 174418 286164
rect 383654 286152 383660 286164
rect 383712 286152 383718 286204
rect 176194 286084 176200 286136
rect 176252 286124 176258 286136
rect 387794 286124 387800 286136
rect 176252 286096 387800 286124
rect 176252 286084 176258 286096
rect 387794 286084 387800 286096
rect 387852 286084 387858 286136
rect 181346 286016 181352 286068
rect 181404 286056 181410 286068
rect 402974 286056 402980 286068
rect 181404 286028 402980 286056
rect 181404 286016 181410 286028
rect 402974 286016 402980 286028
rect 403032 286016 403038 286068
rect 182450 285948 182456 286000
rect 182508 285988 182514 286000
rect 404354 285988 404360 286000
rect 182508 285960 404360 285988
rect 182508 285948 182514 285960
rect 404354 285948 404360 285960
rect 404412 285948 404418 286000
rect 182818 285880 182824 285932
rect 182876 285920 182882 285932
rect 407114 285920 407120 285932
rect 182876 285892 407120 285920
rect 182876 285880 182882 285892
rect 407114 285880 407120 285892
rect 407172 285880 407178 285932
rect 184290 285812 184296 285864
rect 184348 285852 184354 285864
rect 412634 285852 412640 285864
rect 184348 285824 412640 285852
rect 184348 285812 184354 285824
rect 412634 285812 412640 285824
rect 412692 285812 412698 285864
rect 185762 285744 185768 285796
rect 185820 285784 185826 285796
rect 416774 285784 416780 285796
rect 185820 285756 416780 285784
rect 185820 285744 185826 285756
rect 416774 285744 416780 285756
rect 416832 285744 416838 285796
rect 187234 285676 187240 285728
rect 187292 285716 187298 285728
rect 422294 285716 422300 285728
rect 187292 285688 422300 285716
rect 187292 285676 187298 285688
rect 422294 285676 422300 285688
rect 422352 285676 422358 285728
rect 145650 285268 145656 285320
rect 145708 285308 145714 285320
rect 177390 285308 177396 285320
rect 145708 285280 177396 285308
rect 145708 285268 145714 285280
rect 177390 285268 177396 285280
rect 177448 285268 177454 285320
rect 144546 285200 144552 285252
rect 144604 285240 144610 285252
rect 177298 285240 177304 285252
rect 144604 285212 177304 285240
rect 144604 285200 144610 285212
rect 177298 285200 177304 285212
rect 177356 285200 177362 285252
rect 203518 285200 203524 285252
rect 203576 285240 203582 285252
rect 222470 285240 222476 285252
rect 203576 285212 222476 285240
rect 203576 285200 203582 285212
rect 222470 285200 222476 285212
rect 222528 285200 222534 285252
rect 229922 285200 229928 285252
rect 229980 285240 229986 285252
rect 247126 285240 247132 285252
rect 229980 285212 247132 285240
rect 229980 285200 229986 285212
rect 247126 285200 247132 285212
rect 247184 285200 247190 285252
rect 134978 285132 134984 285184
rect 135036 285172 135042 285184
rect 188430 285172 188436 285184
rect 135036 285144 188436 285172
rect 135036 285132 135042 285144
rect 188430 285132 188436 285144
rect 188488 285132 188494 285184
rect 206370 285132 206376 285184
rect 206428 285172 206434 285184
rect 230566 285172 230572 285184
rect 206428 285144 230572 285172
rect 206428 285132 206434 285144
rect 230566 285132 230572 285144
rect 230624 285132 230630 285184
rect 260098 285132 260104 285184
rect 260156 285172 260162 285184
rect 268470 285172 268476 285184
rect 260156 285144 268476 285172
rect 260156 285132 260162 285144
rect 268470 285132 268476 285144
rect 268528 285132 268534 285184
rect 170306 285064 170312 285116
rect 170364 285104 170370 285116
rect 371234 285104 371240 285116
rect 170364 285076 371240 285104
rect 170364 285064 170370 285076
rect 371234 285064 371240 285076
rect 371292 285064 371298 285116
rect 40034 284996 40040 285048
rect 40092 285036 40098 285048
rect 149054 285036 149060 285048
rect 40092 285008 149060 285036
rect 40092 284996 40098 285008
rect 149054 284996 149060 285008
rect 149112 284996 149118 285048
rect 172146 284996 172152 285048
rect 172204 285036 172210 285048
rect 376754 285036 376760 285048
rect 172204 285008 376760 285036
rect 172204 284996 172210 285008
rect 376754 284996 376760 285008
rect 376812 284996 376818 285048
rect 18598 284928 18604 284980
rect 18656 284968 18662 284980
rect 149974 284968 149980 284980
rect 18656 284940 149980 284968
rect 18656 284928 18662 284940
rect 149974 284928 149980 284940
rect 150032 284928 150038 284980
rect 175826 284928 175832 284980
rect 175884 284968 175890 284980
rect 386414 284968 386420 284980
rect 175884 284940 386420 284968
rect 175884 284928 175890 284940
rect 386414 284928 386420 284940
rect 386472 284928 386478 284980
rect 179230 284860 179236 284912
rect 179288 284900 179294 284912
rect 396074 284900 396080 284912
rect 179288 284872 396080 284900
rect 179288 284860 179294 284872
rect 396074 284860 396080 284872
rect 396132 284860 396138 284912
rect 179874 284792 179880 284844
rect 179932 284832 179938 284844
rect 397454 284832 397460 284844
rect 179932 284804 397460 284832
rect 179932 284792 179938 284804
rect 397454 284792 397460 284804
rect 397512 284792 397518 284844
rect 185394 284724 185400 284776
rect 185452 284764 185458 284776
rect 414014 284764 414020 284776
rect 185452 284736 414020 284764
rect 185452 284724 185458 284736
rect 414014 284724 414020 284736
rect 414072 284724 414078 284776
rect 186866 284656 186872 284708
rect 186924 284696 186930 284708
rect 419534 284696 419540 284708
rect 186924 284668 419540 284696
rect 186924 284656 186930 284668
rect 419534 284656 419540 284668
rect 419592 284656 419598 284708
rect 188338 284588 188344 284640
rect 188396 284628 188402 284640
rect 423674 284628 423680 284640
rect 188396 284600 423680 284628
rect 188396 284588 188402 284600
rect 423674 284588 423680 284600
rect 423732 284588 423738 284640
rect 189442 284520 189448 284572
rect 189500 284560 189506 284572
rect 426434 284560 426440 284572
rect 189500 284532 426440 284560
rect 189500 284520 189506 284532
rect 426434 284520 426440 284532
rect 426492 284520 426498 284572
rect 190270 284452 190276 284504
rect 190328 284492 190334 284504
rect 429194 284492 429200 284504
rect 190328 284464 429200 284492
rect 190328 284452 190334 284464
rect 429194 284452 429200 284464
rect 429252 284452 429258 284504
rect 169662 284384 169668 284436
rect 169720 284424 169726 284436
rect 436094 284424 436100 284436
rect 169720 284396 436100 284424
rect 169720 284384 169726 284396
rect 436094 284384 436100 284396
rect 436152 284384 436158 284436
rect 179138 284316 179144 284368
rect 179196 284356 179202 284368
rect 448514 284356 448520 284368
rect 179196 284328 448520 284356
rect 179196 284316 179202 284328
rect 448514 284316 448520 284328
rect 448572 284316 448578 284368
rect 130562 283772 130568 283824
rect 130620 283812 130626 283824
rect 321094 283812 321100 283824
rect 130620 283784 321100 283812
rect 130620 283772 130626 283784
rect 321094 283772 321100 283784
rect 321152 283772 321158 283824
rect 178310 283704 178316 283756
rect 178368 283744 178374 283756
rect 380894 283744 380900 283756
rect 178368 283716 380900 283744
rect 178368 283704 178374 283716
rect 380894 283704 380900 283716
rect 380952 283704 380958 283756
rect 187786 283636 187792 283688
rect 187844 283676 187850 283688
rect 393314 283676 393320 283688
rect 187844 283648 393320 283676
rect 187844 283636 187850 283648
rect 393314 283636 393320 283648
rect 393372 283636 393378 283688
rect 136082 283568 136088 283620
rect 136140 283608 136146 283620
rect 537570 283608 537576 283620
rect 136140 283580 537576 283608
rect 136140 283568 136146 283580
rect 537570 283568 537576 283580
rect 537628 283568 537634 283620
rect 169754 283500 169760 283552
rect 169812 283540 169818 283552
rect 433334 283540 433340 283552
rect 169812 283512 433340 283540
rect 169812 283500 169818 283512
rect 433334 283500 433340 283512
rect 433392 283500 433398 283552
rect 116670 283432 116676 283484
rect 116728 283472 116734 283484
rect 161014 283472 161020 283484
rect 116728 283444 161020 283472
rect 116728 283432 116734 283444
rect 161014 283432 161020 283444
rect 161072 283432 161078 283484
rect 174906 283432 174912 283484
rect 174964 283472 174970 283484
rect 580534 283472 580540 283484
rect 174964 283444 580540 283472
rect 174964 283432 174970 283444
rect 580534 283432 580540 283444
rect 580592 283432 580598 283484
rect 119522 283364 119528 283416
rect 119580 283404 119586 283416
rect 160094 283404 160100 283416
rect 119580 283376 160100 283404
rect 119580 283364 119586 283376
rect 160094 283364 160100 283376
rect 160152 283364 160158 283416
rect 173802 283364 173808 283416
rect 173860 283404 173866 283416
rect 580718 283404 580724 283416
rect 173860 283376 580724 283404
rect 173860 283364 173866 283376
rect 580718 283364 580724 283376
rect 580776 283364 580782 283416
rect 126146 283296 126152 283348
rect 126204 283336 126210 283348
rect 538950 283336 538956 283348
rect 126204 283308 538956 283336
rect 126204 283296 126210 283308
rect 538950 283296 538956 283308
rect 539008 283296 539014 283348
rect 127250 283228 127256 283280
rect 127308 283268 127314 283280
rect 540238 283268 540244 283280
rect 127308 283240 540244 283268
rect 127308 283228 127314 283240
rect 540238 283228 540244 283240
rect 540296 283228 540302 283280
rect 125410 283160 125416 283212
rect 125468 283200 125474 283212
rect 538858 283200 538864 283212
rect 125468 283172 538864 283200
rect 125468 283160 125474 283172
rect 538858 283160 538864 283172
rect 538916 283160 538922 283212
rect 128262 283092 128268 283144
rect 128320 283132 128326 283144
rect 543090 283132 543096 283144
rect 128320 283104 543096 283132
rect 128320 283092 128326 283104
rect 543090 283092 543096 283104
rect 543148 283092 543154 283144
rect 129458 283024 129464 283076
rect 129516 283064 129522 283076
rect 544378 283064 544384 283076
rect 129516 283036 544384 283064
rect 129516 283024 129522 283036
rect 544378 283024 544384 283036
rect 544436 283024 544442 283076
rect 126514 282956 126520 283008
rect 126572 282996 126578 283008
rect 542998 282996 543004 283008
rect 126572 282968 543004 282996
rect 126572 282956 126578 282968
rect 542998 282956 543004 282968
rect 543056 282956 543062 283008
rect 143442 282888 143448 282940
rect 143500 282928 143506 282940
rect 580350 282928 580356 282940
rect 143500 282900 580356 282928
rect 143500 282888 143506 282900
rect 580350 282888 580356 282900
rect 580408 282888 580414 282940
rect 192018 282820 192024 282872
rect 192076 282860 192082 282872
rect 192294 282860 192300 282872
rect 192076 282832 192300 282860
rect 192076 282820 192082 282832
rect 192294 282820 192300 282832
rect 192352 282820 192358 282872
rect 200114 282820 200120 282872
rect 200172 282860 200178 282872
rect 200758 282860 200764 282872
rect 200172 282832 200764 282860
rect 200172 282820 200178 282832
rect 200758 282820 200764 282832
rect 200816 282820 200822 282872
rect 202966 282820 202972 282872
rect 203024 282860 203030 282872
rect 203334 282860 203340 282872
rect 203024 282832 203340 282860
rect 203024 282820 203030 282832
rect 203334 282820 203340 282832
rect 203392 282820 203398 282872
rect 206002 282820 206008 282872
rect 206060 282860 206066 282872
rect 206278 282860 206284 282872
rect 206060 282832 206284 282860
rect 206060 282820 206066 282832
rect 206278 282820 206284 282832
rect 206336 282820 206342 282872
rect 208578 282820 208584 282872
rect 208636 282860 208642 282872
rect 208854 282860 208860 282872
rect 208636 282832 208860 282860
rect 208636 282820 208642 282832
rect 208854 282820 208860 282832
rect 208912 282820 208918 282872
rect 212534 282820 212540 282872
rect 212592 282860 212598 282872
rect 213270 282860 213276 282872
rect 212592 282832 213276 282860
rect 212592 282820 212598 282832
rect 213270 282820 213276 282832
rect 213328 282820 213334 282872
rect 219894 282820 219900 282872
rect 219952 282860 219958 282872
rect 222194 282860 222200 282872
rect 219952 282832 222200 282860
rect 219952 282820 219958 282832
rect 222194 282820 222200 282832
rect 222252 282820 222258 282872
rect 258258 282820 258264 282872
rect 258316 282860 258322 282872
rect 258534 282860 258540 282872
rect 258316 282832 258540 282860
rect 258316 282820 258322 282832
rect 258534 282820 258540 282832
rect 258592 282820 258598 282872
rect 259730 282820 259736 282872
rect 259788 282860 259794 282872
rect 260006 282860 260012 282872
rect 259788 282832 260012 282860
rect 259788 282820 259794 282832
rect 260006 282820 260012 282832
rect 260064 282820 260070 282872
rect 266630 282820 266636 282872
rect 266688 282860 266694 282872
rect 266998 282860 267004 282872
rect 266688 282832 267004 282860
rect 266688 282820 266694 282832
rect 266998 282820 267004 282832
rect 267056 282820 267062 282872
rect 203058 282752 203064 282804
rect 203116 282792 203122 282804
rect 203702 282792 203708 282804
rect 203116 282764 203708 282792
rect 203116 282752 203122 282764
rect 203702 282752 203708 282764
rect 203760 282752 203766 282804
rect 166258 282548 166264 282600
rect 166316 282588 166322 282600
rect 178034 282588 178040 282600
rect 166316 282560 178040 282588
rect 166316 282548 166322 282560
rect 178034 282548 178040 282560
rect 178092 282548 178098 282600
rect 90358 282480 90364 282532
rect 90416 282520 90422 282532
rect 162854 282520 162860 282532
rect 90416 282492 162860 282520
rect 90416 282480 90422 282492
rect 162854 282480 162860 282492
rect 162912 282480 162918 282532
rect 173710 282480 173716 282532
rect 173768 282520 173774 282532
rect 178310 282520 178316 282532
rect 173768 282492 178316 282520
rect 173768 282480 173774 282492
rect 178310 282480 178316 282492
rect 178368 282480 178374 282532
rect 148962 282412 148968 282464
rect 149020 282452 149026 282464
rect 176654 282452 176660 282464
rect 149020 282424 176660 282452
rect 149020 282412 149026 282424
rect 176654 282412 176660 282424
rect 176712 282412 176718 282464
rect 177942 282412 177948 282464
rect 178000 282452 178006 282464
rect 187786 282452 187792 282464
rect 178000 282424 187792 282452
rect 178000 282412 178006 282424
rect 187786 282412 187792 282424
rect 187844 282412 187850 282464
rect 148226 282344 148232 282396
rect 148284 282384 148290 282396
rect 178218 282384 178224 282396
rect 148284 282356 178224 282384
rect 148284 282344 148290 282356
rect 178218 282344 178224 282356
rect 178276 282344 178282 282396
rect 180242 282344 180248 282396
rect 180300 282384 180306 282396
rect 187878 282384 187884 282396
rect 180300 282356 187884 282384
rect 180300 282344 180306 282356
rect 187878 282344 187884 282356
rect 187936 282344 187942 282396
rect 206370 282344 206376 282396
rect 206428 282384 206434 282396
rect 226518 282384 226524 282396
rect 206428 282356 226524 282384
rect 206428 282344 206434 282356
rect 226518 282344 226524 282356
rect 226576 282344 226582 282396
rect 127618 282276 127624 282328
rect 127676 282316 127682 282328
rect 143442 282316 143448 282328
rect 127676 282288 143448 282316
rect 127676 282276 127682 282288
rect 143442 282276 143448 282288
rect 143500 282276 143506 282328
rect 147490 282276 147496 282328
rect 147548 282316 147554 282328
rect 178126 282316 178132 282328
rect 147548 282288 178132 282316
rect 147548 282276 147554 282288
rect 178126 282276 178132 282288
rect 178184 282276 178190 282328
rect 186130 282276 186136 282328
rect 186188 282316 186194 282328
rect 191650 282316 191656 282328
rect 186188 282288 191656 282316
rect 186188 282276 186194 282288
rect 191650 282276 191656 282288
rect 191708 282276 191714 282328
rect 214650 282276 214656 282328
rect 214708 282316 214714 282328
rect 252278 282316 252284 282328
rect 214708 282288 252284 282316
rect 214708 282276 214714 282288
rect 252278 282276 252284 282288
rect 252336 282276 252342 282328
rect 130194 282208 130200 282260
rect 130252 282248 130258 282260
rect 173802 282248 173808 282260
rect 130252 282220 173808 282248
rect 130252 282208 130258 282220
rect 173802 282208 173808 282220
rect 173860 282208 173866 282260
rect 181714 282208 181720 282260
rect 181772 282248 181778 282260
rect 319898 282248 319904 282260
rect 181772 282220 319904 282248
rect 181772 282208 181778 282220
rect 319898 282208 319904 282220
rect 319956 282208 319962 282260
rect 129090 282140 129096 282192
rect 129148 282180 129154 282192
rect 174906 282180 174912 282192
rect 129148 282152 174912 282180
rect 129148 282140 129154 282152
rect 174906 282140 174912 282152
rect 174964 282140 174970 282192
rect 178402 282140 178408 282192
rect 178460 282180 178466 282192
rect 320082 282180 320088 282192
rect 178460 282152 320088 282180
rect 178460 282140 178466 282152
rect 320082 282140 320088 282152
rect 320140 282140 320146 282192
rect 15838 282072 15844 282124
rect 15896 282112 15902 282124
rect 165062 282112 165068 282124
rect 15896 282084 165068 282112
rect 15896 282072 15902 282084
rect 165062 282072 165068 282084
rect 165120 282072 165126 282124
rect 174998 282072 175004 282124
rect 175056 282112 175062 282124
rect 318150 282112 318156 282124
rect 175056 282084 318156 282112
rect 175056 282072 175062 282084
rect 318150 282072 318156 282084
rect 318208 282072 318214 282124
rect 133782 282004 133788 282056
rect 133840 282044 133846 282056
rect 163958 282044 163964 282056
rect 133840 282016 163964 282044
rect 133840 282004 133846 282016
rect 163958 282004 163964 282016
rect 164016 282004 164022 282056
rect 169570 282004 169576 282056
rect 169628 282044 169634 282056
rect 314838 282044 314844 282056
rect 169628 282016 314844 282044
rect 169628 282004 169634 282016
rect 314838 282004 314844 282016
rect 314896 282004 314902 282056
rect 120902 281936 120908 281988
rect 120960 281976 120966 281988
rect 158898 281976 158904 281988
rect 120960 281948 158904 281976
rect 120960 281936 120966 281948
rect 158898 281936 158904 281948
rect 158956 281936 158962 281988
rect 171410 281936 171416 281988
rect 171468 281976 171474 281988
rect 319438 281976 319444 281988
rect 171468 281948 319444 281976
rect 171468 281936 171474 281948
rect 319438 281936 319444 281948
rect 319496 281936 319502 281988
rect 119614 281868 119620 281920
rect 119672 281908 119678 281920
rect 119672 281880 156368 281908
rect 119672 281868 119678 281880
rect 119430 281800 119436 281852
rect 119488 281840 119494 281852
rect 156230 281840 156236 281852
rect 119488 281812 156236 281840
rect 119488 281800 119494 281812
rect 156230 281800 156236 281812
rect 156288 281800 156294 281852
rect 156340 281840 156368 281880
rect 158806 281868 158812 281920
rect 158864 281908 158870 281920
rect 164326 281908 164332 281920
rect 158864 281880 164332 281908
rect 158864 281868 158870 281880
rect 164326 281868 164332 281880
rect 164384 281868 164390 281920
rect 170950 281868 170956 281920
rect 171008 281908 171014 281920
rect 320910 281908 320916 281920
rect 171008 281880 320916 281908
rect 171008 281868 171014 281880
rect 320910 281868 320916 281880
rect 320968 281868 320974 281920
rect 159174 281840 159180 281852
rect 156340 281812 159180 281840
rect 159174 281800 159180 281812
rect 159232 281800 159238 281852
rect 169202 281800 169208 281852
rect 169260 281840 169266 281852
rect 321002 281840 321008 281852
rect 169260 281812 321008 281840
rect 169260 281800 169266 281812
rect 321002 281800 321008 281812
rect 321060 281800 321066 281852
rect 120810 281732 120816 281784
rect 120868 281772 120874 281784
rect 162118 281772 162124 281784
rect 120868 281744 162124 281772
rect 120868 281732 120874 281744
rect 162118 281732 162124 281744
rect 162176 281732 162182 281784
rect 174722 281732 174728 281784
rect 174780 281772 174786 281784
rect 459554 281772 459560 281784
rect 174780 281744 459560 281772
rect 174780 281732 174786 281744
rect 459554 281732 459560 281744
rect 459612 281732 459618 281784
rect 120718 281664 120724 281716
rect 120776 281704 120782 281716
rect 164694 281704 164700 281716
rect 120776 281676 164700 281704
rect 120776 281664 120782 281676
rect 164694 281664 164700 281676
rect 164752 281664 164758 281716
rect 167730 281664 167736 281716
rect 167788 281704 167794 281716
rect 453298 281704 453304 281716
rect 167788 281676 453304 281704
rect 167788 281664 167794 281676
rect 453298 281664 453304 281676
rect 453356 281664 453362 281716
rect 121270 281596 121276 281648
rect 121328 281636 121334 281648
rect 124582 281636 124588 281648
rect 121328 281608 124588 281636
rect 121328 281596 121334 281608
rect 124582 281596 124588 281608
rect 124640 281596 124646 281648
rect 156230 281596 156236 281648
rect 156288 281636 156294 281648
rect 160278 281636 160284 281648
rect 156288 281608 160284 281636
rect 156288 281596 156294 281608
rect 160278 281596 160284 281608
rect 160336 281596 160342 281648
rect 168098 281596 168104 281648
rect 168156 281636 168162 281648
rect 169754 281636 169760 281648
rect 168156 281608 169760 281636
rect 168156 281596 168162 281608
rect 169754 281596 169760 281608
rect 169812 281596 169818 281648
rect 176562 281596 176568 281648
rect 176620 281636 176626 281648
rect 462314 281636 462320 281648
rect 176620 281608 462320 281636
rect 176620 281596 176626 281608
rect 462314 281596 462320 281608
rect 462372 281596 462378 281648
rect 143442 281528 143448 281580
rect 143500 281568 143506 281580
rect 160646 281568 160652 281580
rect 143500 281540 160652 281568
rect 143500 281528 143506 281540
rect 160646 281528 160652 281540
rect 160704 281528 160710 281580
rect 166626 281528 166632 281580
rect 166684 281568 166690 281580
rect 179414 281568 179420 281580
rect 166684 281540 179420 281568
rect 166684 281528 166690 281540
rect 179414 281528 179420 281540
rect 179472 281528 179478 281580
rect 188706 281528 188712 281580
rect 188764 281568 188770 281580
rect 481634 281568 481640 281580
rect 188764 281540 481640 281568
rect 188764 281528 188770 281540
rect 481634 281528 481640 281540
rect 481692 281528 481698 281580
rect 184750 281052 184756 281104
rect 184808 281092 184814 281104
rect 318058 281092 318064 281104
rect 184808 281064 318064 281092
rect 184808 281052 184814 281064
rect 318058 281052 318064 281064
rect 318116 281052 318122 281104
rect 130930 280984 130936 281036
rect 130988 281024 130994 281036
rect 318242 281024 318248 281036
rect 130988 280996 318248 281024
rect 130988 280984 130994 280996
rect 318242 280984 318248 280996
rect 318300 280984 318306 281036
rect 3510 280916 3516 280968
rect 3568 280956 3574 280968
rect 133782 280956 133788 280968
rect 3568 280928 133788 280956
rect 3568 280916 3574 280928
rect 133782 280916 133788 280928
rect 133840 280916 133846 280968
rect 178034 280916 178040 280968
rect 178092 280956 178098 280968
rect 431954 280956 431960 280968
rect 178092 280928 431960 280956
rect 178092 280916 178098 280928
rect 431954 280916 431960 280928
rect 432012 280916 432018 280968
rect 3786 280848 3792 280900
rect 3844 280888 3850 280900
rect 143442 280888 143448 280900
rect 3844 280860 143448 280888
rect 3844 280848 3850 280860
rect 143442 280848 143448 280860
rect 143500 280848 143506 280900
rect 191650 280848 191656 280900
rect 191708 280888 191714 280900
rect 476114 280888 476120 280900
rect 191708 280860 476120 280888
rect 191708 280848 191714 280860
rect 476114 280848 476120 280860
rect 476172 280848 476178 280900
rect 3694 280780 3700 280832
rect 3752 280820 3758 280832
rect 162486 280820 162492 280832
rect 3752 280792 162492 280820
rect 3752 280780 3758 280792
rect 162486 280780 162492 280792
rect 162544 280780 162550 280832
rect 175090 280780 175096 280832
rect 175148 280820 175154 280832
rect 185486 280820 185492 280832
rect 175148 280792 185492 280820
rect 175148 280780 175154 280792
rect 185486 280780 185492 280792
rect 185544 280780 185550 280832
rect 185578 280780 185584 280832
rect 185636 280820 185642 280832
rect 580626 280820 580632 280832
rect 185636 280792 580632 280820
rect 185636 280780 185642 280792
rect 580626 280780 580632 280792
rect 580684 280780 580690 280832
rect 131022 280712 131028 280764
rect 131080 280752 131086 280764
rect 321186 280752 321192 280764
rect 131080 280724 321192 280752
rect 131080 280712 131086 280724
rect 321186 280712 321192 280724
rect 321244 280712 321250 280764
rect 129550 280644 129556 280696
rect 129608 280684 129614 280696
rect 319990 280684 319996 280696
rect 129608 280656 319996 280684
rect 129608 280644 129614 280656
rect 319990 280644 319996 280656
rect 320048 280644 320054 280696
rect 168190 280576 168196 280628
rect 168248 280616 168254 280628
rect 367094 280616 367100 280628
rect 168248 280588 367100 280616
rect 168248 280576 168254 280588
rect 367094 280576 367100 280588
rect 367152 280576 367158 280628
rect 180702 280508 180708 280560
rect 180760 280548 180766 280560
rect 400214 280548 400220 280560
rect 180760 280520 400220 280548
rect 180760 280508 180766 280520
rect 400214 280508 400220 280520
rect 400272 280508 400278 280560
rect 115290 280440 115296 280492
rect 115348 280480 115354 280492
rect 159542 280480 159548 280492
rect 115348 280452 159548 280480
rect 115348 280440 115354 280452
rect 159542 280440 159548 280452
rect 159600 280440 159606 280492
rect 173618 280440 173624 280492
rect 173676 280480 173682 280492
rect 440234 280480 440240 280492
rect 173676 280452 440240 280480
rect 173676 280440 173682 280452
rect 440234 280440 440240 280452
rect 440292 280440 440298 280492
rect 119338 280372 119344 280424
rect 119396 280412 119402 280424
rect 163590 280412 163596 280424
rect 119396 280384 163596 280412
rect 119396 280372 119402 280384
rect 163590 280372 163596 280384
rect 163648 280372 163654 280424
rect 171778 280372 171784 280424
rect 171836 280412 171842 280424
rect 438854 280412 438860 280424
rect 171836 280384 438860 280412
rect 171836 280372 171842 280384
rect 438854 280372 438860 280384
rect 438912 280372 438918 280424
rect 116578 280304 116584 280356
rect 116636 280344 116642 280356
rect 161566 280344 161572 280356
rect 116636 280316 161572 280344
rect 116636 280304 116642 280316
rect 161566 280304 161572 280316
rect 161624 280304 161630 280356
rect 177298 280304 177304 280356
rect 177356 280344 177362 280356
rect 177356 280316 180794 280344
rect 177356 280304 177362 280316
rect 115198 280236 115204 280288
rect 115256 280276 115262 280288
rect 161750 280276 161756 280288
rect 115256 280248 161756 280276
rect 115256 280236 115262 280248
rect 161750 280236 161756 280248
rect 161808 280236 161814 280288
rect 180766 280276 180794 280316
rect 185486 280304 185492 280356
rect 185544 280344 185550 280356
rect 442994 280344 443000 280356
rect 185544 280316 443000 280344
rect 185544 280304 185550 280316
rect 442994 280304 443000 280316
rect 443052 280304 443058 280356
rect 445754 280276 445760 280288
rect 180766 280248 445760 280276
rect 445754 280236 445760 280248
rect 445812 280236 445818 280288
rect 3602 280168 3608 280220
rect 3660 280208 3666 280220
rect 163452 280208 163458 280220
rect 3660 280180 163458 280208
rect 3660 280168 3666 280180
rect 163452 280168 163458 280180
rect 163510 280168 163516 280220
rect 165660 280168 165666 280220
rect 165718 280208 165724 280220
rect 511258 280208 511264 280220
rect 165718 280180 511264 280208
rect 165718 280168 165724 280180
rect 511258 280168 511264 280180
rect 511316 280168 511322 280220
rect 121362 280100 121368 280152
rect 121420 280140 121426 280152
rect 124214 280140 124220 280152
rect 121420 280112 124220 280140
rect 121420 280100 121426 280112
rect 124214 280100 124220 280112
rect 124272 280100 124278 280152
rect 314838 279828 314844 279880
rect 314896 279868 314902 279880
rect 491294 279868 491300 279880
rect 314896 279840 491300 279868
rect 314896 279828 314902 279840
rect 491294 279828 491300 279840
rect 491352 279828 491358 279880
rect 179414 279760 179420 279812
rect 179472 279800 179478 279812
rect 361666 279800 361672 279812
rect 179472 279772 361672 279800
rect 179472 279760 179478 279772
rect 361666 279760 361672 279772
rect 361724 279760 361730 279812
rect 187878 279692 187884 279744
rect 187936 279732 187942 279744
rect 467834 279732 467840 279744
rect 187936 279704 467840 279732
rect 187936 279692 187942 279704
rect 467834 279692 467840 279704
rect 467892 279692 467898 279744
rect 177666 279624 177672 279676
rect 177724 279664 177730 279676
rect 390554 279664 390560 279676
rect 177724 279636 390560 279664
rect 177724 279624 177730 279636
rect 390554 279624 390560 279636
rect 390612 279624 390618 279676
rect 158806 279596 158812 279608
rect 142126 279568 158812 279596
rect 3418 279488 3424 279540
rect 3476 279528 3482 279540
rect 142126 279528 142154 279568
rect 158806 279556 158812 279568
rect 158864 279556 158870 279608
rect 180610 279556 180616 279608
rect 180668 279596 180674 279608
rect 180668 279568 180794 279596
rect 180668 279556 180674 279568
rect 3476 279500 142154 279528
rect 180766 279528 180794 279568
rect 183922 279556 183928 279608
rect 183980 279596 183986 279608
rect 409874 279596 409880 279608
rect 183980 279568 409880 279596
rect 183980 279556 183986 279568
rect 409874 279556 409880 279568
rect 409932 279556 409938 279608
rect 505094 279528 505100 279540
rect 180766 279500 505100 279528
rect 3476 279488 3482 279500
rect 505094 279488 505100 279500
rect 505152 279488 505158 279540
rect 3326 267656 3332 267708
rect 3384 267696 3390 267708
rect 120902 267696 120908 267708
rect 3384 267668 120908 267696
rect 3384 267656 3390 267668
rect 120902 267656 120908 267668
rect 120960 267656 120966 267708
rect 321186 259360 321192 259412
rect 321244 259400 321250 259412
rect 579798 259400 579804 259412
rect 321244 259372 579804 259400
rect 321244 259360 321250 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 2958 255212 2964 255264
rect 3016 255252 3022 255264
rect 115290 255252 115296 255264
rect 3016 255224 115296 255252
rect 3016 255212 3022 255224
rect 115290 255212 115296 255224
rect 115348 255212 115354 255264
rect 321094 245556 321100 245608
rect 321152 245596 321158 245608
rect 580166 245596 580172 245608
rect 321152 245568 580172 245596
rect 321152 245556 321158 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3326 241408 3332 241460
rect 3384 241448 3390 241460
rect 119614 241448 119620 241460
rect 3384 241420 119620 241448
rect 3384 241408 3390 241420
rect 119614 241408 119620 241420
rect 119672 241408 119678 241460
rect 320082 233928 320088 233980
rect 320140 233968 320146 233980
rect 465442 233968 465448 233980
rect 320140 233940 465448 233968
rect 320140 233928 320146 233940
rect 465442 233928 465448 233940
rect 465500 233928 465506 233980
rect 319438 233860 319444 233912
rect 319496 233900 319502 233912
rect 494146 233900 494152 233912
rect 319496 233872 494152 233900
rect 319496 233860 319502 233872
rect 494146 233860 494152 233872
rect 494204 233860 494210 233912
rect 319990 233180 319996 233232
rect 320048 233220 320054 233232
rect 579982 233220 579988 233232
rect 320048 233192 579988 233220
rect 320048 233180 320054 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 321002 232976 321008 233028
rect 321060 233016 321066 233028
rect 453206 233016 453212 233028
rect 321060 232988 453212 233016
rect 321060 232976 321066 232988
rect 453206 232976 453212 232988
rect 453264 232976 453270 233028
rect 453298 232976 453304 233028
rect 453356 233016 453362 233028
rect 489362 233016 489368 233028
rect 453356 232988 489368 233016
rect 453356 232976 453362 232988
rect 489362 232976 489368 232988
rect 489420 232976 489426 233028
rect 491938 232976 491944 233028
rect 491996 233016 492002 233028
rect 503714 233016 503720 233028
rect 491996 232988 503720 233016
rect 491996 232976 492002 232988
rect 503714 232976 503720 232988
rect 503772 232976 503778 233028
rect 320910 232908 320916 232960
rect 320968 232948 320974 232960
rect 455874 232948 455880 232960
rect 320968 232920 455880 232948
rect 320968 232908 320974 232920
rect 455874 232908 455880 232920
rect 455932 232908 455938 232960
rect 456058 232908 456064 232960
rect 456116 232948 456122 232960
rect 520458 232948 520464 232960
rect 456116 232920 520464 232948
rect 456116 232908 456122 232920
rect 520458 232908 520464 232920
rect 520516 232908 520522 232960
rect 319898 232840 319904 232892
rect 319956 232880 319962 232892
rect 469766 232880 469772 232892
rect 319956 232852 469772 232880
rect 319956 232840 319962 232852
rect 469766 232840 469772 232852
rect 469824 232840 469830 232892
rect 469858 232840 469864 232892
rect 469916 232880 469922 232892
rect 525242 232880 525248 232892
rect 469916 232852 525248 232880
rect 469916 232840 469922 232852
rect 525242 232840 525248 232852
rect 525300 232840 525306 232892
rect 319714 232772 319720 232824
rect 319772 232812 319778 232824
rect 496538 232812 496544 232824
rect 319772 232784 496544 232812
rect 319772 232772 319778 232784
rect 496538 232772 496544 232784
rect 496596 232772 496602 232824
rect 319530 232704 319536 232756
rect 319588 232744 319594 232756
rect 501322 232744 501328 232756
rect 319588 232716 501328 232744
rect 319588 232704 319594 232716
rect 501322 232704 501328 232716
rect 501380 232704 501386 232756
rect 320818 232636 320824 232688
rect 320876 232676 320882 232688
rect 508498 232676 508504 232688
rect 320876 232648 508504 232676
rect 320876 232636 320882 232648
rect 508498 232636 508504 232648
rect 508556 232636 508562 232688
rect 319806 232568 319812 232620
rect 319864 232608 319870 232620
rect 510890 232608 510896 232620
rect 319864 232580 510896 232608
rect 319864 232568 319870 232580
rect 510890 232568 510896 232580
rect 510948 232568 510954 232620
rect 511258 232568 511264 232620
rect 511316 232608 511322 232620
rect 527634 232608 527640 232620
rect 511316 232580 527640 232608
rect 511316 232568 511322 232580
rect 527634 232568 527640 232580
rect 527692 232568 527698 232620
rect 319622 232500 319628 232552
rect 319680 232540 319686 232552
rect 522850 232540 522856 232552
rect 319680 232512 522856 232540
rect 319680 232500 319686 232512
rect 522850 232500 522856 232512
rect 522908 232500 522914 232552
rect 319438 231820 319444 231872
rect 319496 231860 319502 231872
rect 537202 231860 537208 231872
rect 319496 231832 537208 231860
rect 319496 231820 319502 231832
rect 537202 231820 537208 231832
rect 537260 231820 537266 231872
rect 319530 230460 319536 230512
rect 319588 230500 319594 230512
rect 530026 230500 530032 230512
rect 319588 230472 530032 230500
rect 319588 230460 319594 230472
rect 530026 230460 530032 230472
rect 530084 230460 530090 230512
rect 3050 215228 3056 215280
rect 3108 215268 3114 215280
rect 119522 215268 119528 215280
rect 3108 215240 119528 215268
rect 3108 215228 3114 215240
rect 119522 215228 119528 215240
rect 119580 215228 119586 215280
rect 544378 206932 544384 206984
rect 544436 206972 544442 206984
rect 580166 206972 580172 206984
rect 544436 206944 580172 206972
rect 544436 206932 544442 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3326 188980 3332 189032
rect 3384 189020 3390 189032
rect 119430 189020 119436 189032
rect 3384 188992 119436 189020
rect 3384 188980 3390 188992
rect 119430 188980 119436 188992
rect 119488 188980 119494 189032
rect 543090 166948 543096 167000
rect 543148 166988 543154 167000
rect 580166 166988 580172 167000
rect 543148 166960 580172 166988
rect 543148 166948 543154 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3050 164160 3056 164212
rect 3108 164200 3114 164212
rect 116670 164200 116676 164212
rect 3108 164172 116676 164200
rect 3108 164160 3114 164172
rect 116670 164160 116676 164172
rect 116728 164160 116734 164212
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 115198 150396 115204 150408
rect 3384 150368 115204 150396
rect 3384 150356 3390 150368
rect 115198 150356 115204 150368
rect 115256 150356 115262 150408
rect 540330 139340 540336 139392
rect 540388 139380 540394 139392
rect 579798 139380 579804 139392
rect 540388 139352 579804 139380
rect 540388 139340 540394 139352
rect 579798 139340 579804 139352
rect 579856 139340 579862 139392
rect 3326 137912 3332 137964
rect 3384 137952 3390 137964
rect 116578 137952 116584 137964
rect 3384 137924 116584 137952
rect 3384 137912 3390 137924
rect 116578 137912 116584 137924
rect 116636 137912 116642 137964
rect 540238 126896 540244 126948
rect 540296 126936 540302 126948
rect 580166 126936 580172 126948
rect 540296 126908 580172 126936
rect 540296 126896 540302 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 542998 113092 543004 113144
rect 543056 113132 543062 113144
rect 579614 113132 579620 113144
rect 543056 113104 579620 113132
rect 543056 113092 543062 113104
rect 579614 113092 579620 113104
rect 579672 113092 579678 113144
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 120810 111772 120816 111784
rect 3384 111744 120816 111772
rect 3384 111732 3390 111744
rect 120810 111732 120816 111744
rect 120868 111732 120874 111784
rect 3326 97928 3332 97980
rect 3384 97968 3390 97980
rect 90358 97968 90364 97980
rect 3384 97940 90364 97968
rect 3384 97928 3390 97940
rect 90358 97928 90364 97940
rect 90416 97928 90422 97980
rect 538950 86912 538956 86964
rect 539008 86952 539014 86964
rect 580166 86952 580172 86964
rect 539008 86924 580172 86952
rect 539008 86912 539014 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 314102 80588 314108 80640
rect 314160 80628 314166 80640
rect 318058 80628 318064 80640
rect 314160 80600 318064 80628
rect 314160 80588 314166 80600
rect 318058 80588 318064 80600
rect 318116 80588 318122 80640
rect 318242 78684 318248 78736
rect 318300 78724 318306 78736
rect 358814 78724 358820 78736
rect 318300 78696 358820 78724
rect 318300 78684 318306 78696
rect 358814 78684 358820 78696
rect 358872 78684 358878 78736
rect 225782 78616 225788 78668
rect 225840 78656 225846 78668
rect 231118 78656 231124 78668
rect 225840 78628 231124 78656
rect 225840 78616 225846 78628
rect 231118 78616 231124 78628
rect 231176 78616 231182 78668
rect 234062 78616 234068 78668
rect 234120 78656 234126 78668
rect 239398 78656 239404 78668
rect 234120 78628 239404 78656
rect 234120 78616 234126 78628
rect 239398 78616 239404 78628
rect 239456 78616 239462 78668
rect 312722 78616 312728 78668
rect 312780 78656 312786 78668
rect 318334 78656 318340 78668
rect 312780 78628 318340 78656
rect 312780 78616 312786 78628
rect 318334 78616 318340 78628
rect 318392 78616 318398 78668
rect 188522 78548 188528 78600
rect 188580 78588 188586 78600
rect 199378 78588 199384 78600
rect 188580 78560 199384 78588
rect 188580 78548 188586 78560
rect 199378 78548 199384 78560
rect 199436 78548 199442 78600
rect 189902 78480 189908 78532
rect 189960 78520 189966 78532
rect 203518 78520 203524 78532
rect 189960 78492 203524 78520
rect 189960 78480 189966 78492
rect 203518 78480 203524 78492
rect 203576 78480 203582 78532
rect 315482 78480 315488 78532
rect 315540 78520 315546 78532
rect 319438 78520 319444 78532
rect 315540 78492 319444 78520
rect 315540 78480 315546 78492
rect 319438 78480 319444 78492
rect 319496 78480 319502 78532
rect 191282 78412 191288 78464
rect 191340 78452 191346 78464
rect 206278 78452 206284 78464
rect 191340 78424 206284 78452
rect 191340 78412 191346 78424
rect 206278 78412 206284 78424
rect 206336 78412 206342 78464
rect 311342 78412 311348 78464
rect 311400 78452 311406 78464
rect 319530 78452 319536 78464
rect 311400 78424 319536 78452
rect 311400 78412 311406 78424
rect 319530 78412 319536 78424
rect 319588 78412 319594 78464
rect 192662 78344 192668 78396
rect 192720 78384 192726 78396
rect 210418 78384 210424 78396
rect 192720 78356 210424 78384
rect 192720 78344 192726 78356
rect 210418 78344 210424 78356
rect 210476 78344 210482 78396
rect 195422 78276 195428 78328
rect 195480 78316 195486 78328
rect 214558 78316 214564 78328
rect 195480 78288 214564 78316
rect 195480 78276 195486 78288
rect 214558 78276 214564 78288
rect 214616 78276 214622 78328
rect 304442 78276 304448 78328
rect 304500 78316 304506 78328
rect 327718 78316 327724 78328
rect 304500 78288 327724 78316
rect 304500 78276 304506 78288
rect 327718 78276 327724 78288
rect 327776 78276 327782 78328
rect 194042 78208 194048 78260
rect 194100 78248 194106 78260
rect 213178 78248 213184 78260
rect 194100 78220 213184 78248
rect 194100 78208 194106 78220
rect 213178 78208 213184 78220
rect 213236 78208 213242 78260
rect 307202 78208 307208 78260
rect 307260 78248 307266 78260
rect 331858 78248 331864 78260
rect 307260 78220 331864 78248
rect 307260 78208 307266 78220
rect 331858 78208 331864 78220
rect 331916 78208 331922 78260
rect 159542 78140 159548 78192
rect 159600 78180 159606 78192
rect 208394 78180 208400 78192
rect 159600 78152 208400 78180
rect 159600 78140 159606 78152
rect 208394 78140 208400 78152
rect 208452 78140 208458 78192
rect 305822 78140 305828 78192
rect 305880 78180 305886 78192
rect 330478 78180 330484 78192
rect 305880 78152 330484 78180
rect 305880 78140 305886 78152
rect 330478 78140 330484 78152
rect 330536 78140 330542 78192
rect 160922 78072 160928 78124
rect 160980 78112 160986 78124
rect 211154 78112 211160 78124
rect 160980 78084 211160 78112
rect 160980 78072 160986 78084
rect 211154 78072 211160 78084
rect 211212 78072 211218 78124
rect 261662 78072 261668 78124
rect 261720 78112 261726 78124
rect 323578 78112 323584 78124
rect 261720 78084 323584 78112
rect 261720 78072 261726 78084
rect 323578 78072 323584 78084
rect 323636 78072 323642 78124
rect 1394 78004 1400 78056
rect 1452 78044 1458 78056
rect 123018 78044 123024 78056
rect 1452 78016 123024 78044
rect 1452 78004 1458 78016
rect 123018 78004 123024 78016
rect 123076 78004 123082 78056
rect 162302 78004 162308 78056
rect 162360 78044 162366 78056
rect 215294 78044 215300 78056
rect 162360 78016 215300 78044
rect 162360 78004 162366 78016
rect 215294 78004 215300 78016
rect 215352 78004 215358 78056
rect 236822 78004 236828 78056
rect 236880 78044 236886 78056
rect 242158 78044 242164 78056
rect 236880 78016 242164 78044
rect 236880 78004 236886 78016
rect 242158 78004 242164 78016
rect 242216 78004 242222 78056
rect 256142 78004 256148 78056
rect 256200 78044 256206 78056
rect 320818 78044 320824 78056
rect 256200 78016 320824 78044
rect 256200 78004 256206 78016
rect 320818 78004 320824 78016
rect 320876 78004 320882 78056
rect 14 77936 20 77988
rect 72 77976 78 77988
rect 121638 77976 121644 77988
rect 72 77948 121644 77976
rect 72 77936 78 77948
rect 121638 77936 121644 77948
rect 121696 77936 121702 77988
rect 163682 77936 163688 77988
rect 163740 77976 163746 77988
rect 218054 77976 218060 77988
rect 163740 77948 218060 77976
rect 163740 77936 163746 77948
rect 218054 77936 218060 77948
rect 218112 77936 218118 77988
rect 218882 77936 218888 77988
rect 218940 77976 218946 77988
rect 228358 77976 228364 77988
rect 218940 77948 228364 77976
rect 218940 77936 218946 77948
rect 228358 77936 228364 77948
rect 228416 77936 228422 77988
rect 247862 77936 247868 77988
rect 247920 77976 247926 77988
rect 313918 77976 313924 77988
rect 247920 77948 313924 77976
rect 247920 77936 247926 77948
rect 313918 77936 313924 77948
rect 313976 77936 313982 77988
rect 239582 77392 239588 77444
rect 239640 77432 239646 77444
rect 244918 77432 244924 77444
rect 239640 77404 244924 77432
rect 239640 77392 239646 77404
rect 244918 77392 244924 77404
rect 244976 77392 244982 77444
rect 242342 77324 242348 77376
rect 242400 77364 242406 77376
rect 246298 77364 246304 77376
rect 242400 77336 246304 77364
rect 242400 77324 242406 77336
rect 246298 77324 246304 77336
rect 246356 77324 246362 77376
rect 125042 77256 125048 77308
rect 125100 77296 125106 77308
rect 125594 77296 125600 77308
rect 125100 77268 125600 77296
rect 125100 77256 125106 77268
rect 125594 77256 125600 77268
rect 125652 77256 125658 77308
rect 129182 77256 129188 77308
rect 129240 77296 129246 77308
rect 129734 77296 129740 77308
rect 129240 77268 129740 77296
rect 129240 77256 129246 77268
rect 129734 77256 129740 77268
rect 129792 77256 129798 77308
rect 155402 77256 155408 77308
rect 155460 77296 155466 77308
rect 156598 77296 156604 77308
rect 155460 77268 156604 77296
rect 155460 77256 155466 77268
rect 156598 77256 156604 77268
rect 156656 77256 156662 77308
rect 156782 77256 156788 77308
rect 156840 77296 156846 77308
rect 157978 77296 157984 77308
rect 156840 77268 157984 77296
rect 156840 77256 156846 77268
rect 157978 77256 157984 77268
rect 158036 77256 158042 77308
rect 158162 77256 158168 77308
rect 158220 77296 158226 77308
rect 159358 77296 159364 77308
rect 158220 77268 159364 77296
rect 158220 77256 158226 77268
rect 159358 77256 159364 77268
rect 159416 77256 159422 77308
rect 171962 77256 171968 77308
rect 172020 77296 172026 77308
rect 173158 77296 173164 77308
rect 172020 77268 173164 77296
rect 172020 77256 172026 77268
rect 173158 77256 173164 77268
rect 173216 77256 173222 77308
rect 214742 77256 214748 77308
rect 214800 77296 214806 77308
rect 217318 77296 217324 77308
rect 214800 77268 217324 77296
rect 214800 77256 214806 77268
rect 217318 77256 217324 77268
rect 217376 77256 217382 77308
rect 221642 77256 221648 77308
rect 221700 77296 221706 77308
rect 224218 77296 224224 77308
rect 221700 77268 224224 77296
rect 221700 77256 221706 77268
rect 224218 77256 224224 77268
rect 224276 77256 224282 77308
rect 240962 77256 240968 77308
rect 241020 77296 241026 77308
rect 242250 77296 242256 77308
rect 241020 77268 242256 77296
rect 241020 77256 241026 77268
rect 242250 77256 242256 77268
rect 242308 77256 242314 77308
rect 245102 77256 245108 77308
rect 245160 77296 245166 77308
rect 247678 77296 247684 77308
rect 245160 77268 247684 77296
rect 245160 77256 245166 77268
rect 247678 77256 247684 77268
rect 247736 77256 247742 77308
rect 165062 75148 165068 75200
rect 165120 75188 165126 75200
rect 222194 75188 222200 75200
rect 165120 75160 222200 75188
rect 165120 75148 165126 75160
rect 222194 75148 222200 75160
rect 222252 75148 222258 75200
rect 195974 73788 195980 73840
rect 196032 73828 196038 73840
rect 303614 73828 303620 73840
rect 196032 73800 303620 73828
rect 196032 73788 196038 73800
rect 303614 73788 303620 73800
rect 303672 73788 303678 73840
rect 538950 73108 538956 73160
rect 539008 73148 539014 73160
rect 579982 73148 579988 73160
rect 539008 73120 579988 73148
rect 539008 73108 539014 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 224218 48968 224224 49020
rect 224276 49008 224282 49020
rect 367094 49008 367100 49020
rect 224276 48980 367100 49008
rect 224276 48968 224282 48980
rect 367094 48968 367100 48980
rect 367152 48968 367158 49020
rect 309134 48220 309140 48272
rect 309192 48260 309198 48272
rect 494882 48260 494888 48272
rect 309192 48232 494888 48260
rect 309192 48220 309198 48232
rect 494882 48220 494888 48232
rect 494940 48220 494946 48272
rect 307754 48152 307760 48204
rect 307812 48192 307818 48204
rect 361574 48192 361580 48204
rect 307812 48164 361580 48192
rect 307812 48152 307818 48164
rect 361574 48152 361580 48164
rect 361632 48192 361638 48204
rect 404906 48192 404912 48204
rect 361632 48164 404912 48192
rect 361632 48152 361638 48164
rect 404906 48152 404912 48164
rect 404964 48152 404970 48204
rect 121270 46860 121276 46912
rect 121328 46900 121334 46912
rect 580166 46900 580172 46912
rect 121328 46872 580172 46900
rect 121328 46860 121334 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 119338 45540 119344 45552
rect 3568 45512 119344 45540
rect 3568 45500 3574 45512
rect 119338 45500 119344 45512
rect 119396 45500 119402 45552
rect 212534 44888 212540 44940
rect 212592 44928 212598 44940
rect 346394 44928 346400 44940
rect 212592 44900 346400 44928
rect 212592 44888 212598 44900
rect 346394 44888 346400 44900
rect 346452 44888 346458 44940
rect 242250 44820 242256 44872
rect 242308 44860 242314 44872
rect 416774 44860 416780 44872
rect 242308 44832 416780 44860
rect 242308 44820 242314 44832
rect 416774 44820 416780 44832
rect 416832 44820 416838 44872
rect 227714 43460 227720 43512
rect 227772 43500 227778 43512
rect 385034 43500 385040 43512
rect 227772 43472 385040 43500
rect 227772 43460 227778 43472
rect 385034 43460 385040 43472
rect 385092 43460 385098 43512
rect 168374 43392 168380 43444
rect 168432 43432 168438 43444
rect 233234 43432 233240 43444
rect 168432 43404 233240 43432
rect 168432 43392 168438 43404
rect 233234 43392 233240 43404
rect 233292 43392 233298 43444
rect 300854 43392 300860 43444
rect 300912 43432 300918 43444
rect 572714 43432 572720 43444
rect 300912 43404 572720 43432
rect 300912 43392 300918 43404
rect 572714 43392 572720 43404
rect 572772 43392 572778 43444
rect 271874 42032 271880 42084
rect 271932 42072 271938 42084
rect 498194 42072 498200 42084
rect 271932 42044 498200 42072
rect 271932 42032 271938 42044
rect 498194 42032 498200 42044
rect 498252 42032 498258 42084
rect 264974 40672 264980 40724
rect 265032 40712 265038 40724
rect 481634 40712 481640 40724
rect 265032 40684 481640 40712
rect 265032 40672 265038 40684
rect 481634 40672 481640 40684
rect 481692 40672 481698 40724
rect 231854 39380 231860 39432
rect 231912 39420 231918 39432
rect 396074 39420 396080 39432
rect 231912 39392 396080 39420
rect 231912 39380 231918 39392
rect 396074 39380 396080 39392
rect 396132 39380 396138 39432
rect 296714 39312 296720 39364
rect 296772 39352 296778 39364
rect 563054 39352 563060 39364
rect 296772 39324 563060 39352
rect 296772 39312 296778 39324
rect 563054 39312 563060 39324
rect 563112 39312 563118 39364
rect 222286 37952 222292 38004
rect 222344 37992 222350 38004
rect 371234 37992 371240 38004
rect 222344 37964 371240 37992
rect 222344 37952 222350 37964
rect 371234 37952 371240 37964
rect 371292 37952 371298 38004
rect 245654 37884 245660 37936
rect 245712 37924 245718 37936
rect 431954 37924 431960 37936
rect 245712 37896 431960 37924
rect 245712 37884 245718 37896
rect 431954 37884 431960 37896
rect 432012 37884 432018 37936
rect 215386 36524 215392 36576
rect 215444 36564 215450 36576
rect 353294 36564 353300 36576
rect 215444 36536 353300 36564
rect 215444 36524 215450 36536
rect 353294 36524 353300 36536
rect 353352 36524 353358 36576
rect 216674 35164 216680 35216
rect 216732 35204 216738 35216
rect 357434 35204 357440 35216
rect 216732 35176 357440 35204
rect 216732 35164 216738 35176
rect 357434 35164 357440 35176
rect 357492 35164 357498 35216
rect 230474 33736 230480 33788
rect 230532 33776 230538 33788
rect 391934 33776 391940 33788
rect 230532 33748 391940 33776
rect 230532 33736 230538 33748
rect 391934 33736 391940 33748
rect 391992 33736 391998 33788
rect 229094 31016 229100 31068
rect 229152 31056 229158 31068
rect 389174 31056 389180 31068
rect 229152 31028 389180 31056
rect 229152 31016 229158 31028
rect 389174 31016 389180 31028
rect 389232 31016 389238 31068
rect 226334 29656 226340 29708
rect 226392 29696 226398 29708
rect 382274 29696 382280 29708
rect 226392 29668 382280 29696
rect 226392 29656 226398 29668
rect 382274 29656 382280 29668
rect 382332 29656 382338 29708
rect 302234 29588 302240 29640
rect 302292 29628 302298 29640
rect 576854 29628 576860 29640
rect 302292 29600 576860 29628
rect 302292 29588 302298 29600
rect 576854 29588 576860 29600
rect 576912 29588 576918 29640
rect 244918 28296 244924 28348
rect 244976 28336 244982 28348
rect 414014 28336 414020 28348
rect 244976 28308 414020 28336
rect 244976 28296 244982 28308
rect 414014 28296 414020 28308
rect 414072 28296 414078 28348
rect 276014 28228 276020 28280
rect 276072 28268 276078 28280
rect 509234 28268 509240 28280
rect 276072 28240 509240 28268
rect 276072 28228 276078 28240
rect 509234 28228 509240 28240
rect 509292 28228 509298 28280
rect 231118 26936 231124 26988
rect 231176 26976 231182 26988
rect 378134 26976 378140 26988
rect 231176 26948 378140 26976
rect 231176 26936 231182 26948
rect 378134 26936 378140 26948
rect 378192 26936 378198 26988
rect 299474 26868 299480 26920
rect 299532 26908 299538 26920
rect 569954 26908 569960 26920
rect 299532 26880 569960 26908
rect 299532 26868 299538 26880
rect 569954 26868 569960 26880
rect 570012 26868 570018 26920
rect 223574 25576 223580 25628
rect 223632 25616 223638 25628
rect 373994 25616 374000 25628
rect 223632 25588 374000 25616
rect 223632 25576 223638 25588
rect 373994 25576 374000 25588
rect 374052 25576 374058 25628
rect 298094 25508 298100 25560
rect 298152 25548 298158 25560
rect 565814 25548 565820 25560
rect 298152 25520 565820 25548
rect 298152 25508 298158 25520
rect 565814 25508 565820 25520
rect 565872 25508 565878 25560
rect 242158 24148 242164 24200
rect 242216 24188 242222 24200
rect 407114 24188 407120 24200
rect 242216 24160 407120 24188
rect 242216 24148 242222 24160
rect 407114 24148 407120 24160
rect 407172 24148 407178 24200
rect 292574 24080 292580 24132
rect 292632 24120 292638 24132
rect 552014 24120 552020 24132
rect 292632 24092 552020 24120
rect 292632 24080 292638 24092
rect 552014 24080 552020 24092
rect 552072 24080 552078 24132
rect 239398 22788 239404 22840
rect 239456 22828 239462 22840
rect 398834 22828 398840 22840
rect 239456 22800 398840 22828
rect 239456 22788 239462 22800
rect 398834 22788 398840 22800
rect 398892 22788 398898 22840
rect 295334 22720 295340 22772
rect 295392 22760 295398 22772
rect 558914 22760 558920 22772
rect 295392 22732 558920 22760
rect 295392 22720 295398 22732
rect 558914 22720 558920 22732
rect 558972 22720 558978 22772
rect 219434 21428 219440 21480
rect 219492 21468 219498 21480
rect 364334 21468 364340 21480
rect 219492 21440 364340 21468
rect 219492 21428 219498 21440
rect 364334 21428 364340 21440
rect 364392 21428 364398 21480
rect 293954 21360 293960 21412
rect 294012 21400 294018 21412
rect 556154 21400 556160 21412
rect 294012 21372 556160 21400
rect 294012 21360 294018 21372
rect 556154 21360 556160 21372
rect 556212 21360 556218 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 15838 20652 15844 20664
rect 3476 20624 15844 20652
rect 3476 20612 3482 20624
rect 15838 20612 15844 20624
rect 15896 20612 15902 20664
rect 121362 20612 121368 20664
rect 121420 20652 121426 20664
rect 579982 20652 579988 20664
rect 121420 20624 579988 20652
rect 121420 20612 121426 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 217318 19932 217324 19984
rect 217376 19972 217382 19984
rect 349154 19972 349160 19984
rect 217376 19944 349160 19972
rect 217376 19932 217382 19944
rect 349154 19932 349160 19944
rect 349212 19932 349218 19984
rect 228358 18640 228364 18692
rect 228416 18680 228422 18692
rect 360194 18680 360200 18692
rect 228416 18652 360200 18680
rect 228416 18640 228422 18652
rect 360194 18640 360200 18652
rect 360252 18640 360258 18692
rect 172514 18572 172520 18624
rect 172572 18612 172578 18624
rect 242986 18612 242992 18624
rect 172572 18584 242992 18612
rect 172572 18572 172578 18584
rect 242986 18572 242992 18584
rect 243044 18572 243050 18624
rect 291194 18572 291200 18624
rect 291252 18612 291258 18624
rect 547874 18612 547880 18624
rect 291252 18584 547880 18612
rect 291252 18572 291258 18584
rect 547874 18572 547880 18584
rect 547932 18572 547938 18624
rect 247678 17280 247684 17332
rect 247736 17320 247742 17332
rect 427814 17320 427820 17332
rect 247736 17292 427820 17320
rect 247736 17280 247742 17292
rect 427814 17280 427820 17292
rect 427872 17280 427878 17332
rect 274634 17212 274640 17264
rect 274692 17252 274698 17264
rect 506474 17252 506480 17264
rect 274692 17224 506480 17252
rect 274692 17212 274698 17224
rect 506474 17212 506480 17224
rect 506532 17212 506538 17264
rect 258074 15920 258080 15972
rect 258132 15960 258138 15972
rect 463970 15960 463976 15972
rect 258132 15932 463976 15960
rect 258132 15920 258138 15932
rect 463970 15920 463976 15932
rect 464028 15920 464034 15972
rect 169754 15852 169760 15904
rect 169812 15892 169818 15904
rect 236546 15892 236552 15904
rect 169812 15864 236552 15892
rect 169812 15852 169818 15864
rect 236546 15852 236552 15864
rect 236604 15852 236610 15904
rect 273254 15852 273260 15904
rect 273312 15892 273318 15904
rect 502978 15892 502984 15904
rect 273312 15864 502984 15892
rect 273312 15852 273318 15864
rect 502978 15852 502984 15864
rect 503036 15852 503042 15904
rect 246298 14492 246304 14544
rect 246356 14532 246362 14544
rect 420914 14532 420920 14544
rect 246356 14504 420920 14532
rect 246356 14492 246362 14504
rect 420914 14492 420920 14504
rect 420972 14492 420978 14544
rect 166994 14424 167000 14476
rect 167052 14464 167058 14476
rect 229370 14464 229376 14476
rect 167052 14436 229376 14464
rect 167052 14424 167058 14436
rect 229370 14424 229376 14436
rect 229428 14424 229434 14476
rect 270494 14424 270500 14476
rect 270552 14464 270558 14476
rect 495434 14464 495440 14476
rect 270552 14436 495440 14464
rect 270552 14424 270558 14436
rect 495434 14424 495440 14436
rect 495492 14424 495498 14476
rect 249794 13132 249800 13184
rect 249852 13172 249858 13184
rect 442626 13172 442632 13184
rect 249852 13144 442632 13172
rect 249852 13132 249858 13144
rect 442626 13132 442632 13144
rect 442684 13132 442690 13184
rect 165614 13064 165620 13116
rect 165672 13104 165678 13116
rect 226334 13104 226340 13116
rect 165672 13076 226340 13104
rect 165672 13064 165678 13076
rect 226334 13064 226340 13076
rect 226392 13064 226398 13116
rect 269114 13064 269120 13116
rect 269172 13104 269178 13116
rect 492306 13104 492312 13116
rect 269172 13076 492312 13104
rect 269172 13064 269178 13076
rect 492306 13064 492312 13076
rect 492364 13064 492370 13116
rect 197354 11772 197360 11824
rect 197412 11812 197418 11824
rect 307938 11812 307944 11824
rect 197412 11784 307944 11812
rect 197412 11772 197418 11784
rect 307938 11772 307944 11784
rect 307996 11772 308002 11824
rect 159358 11704 159364 11756
rect 159416 11744 159422 11756
rect 205082 11744 205088 11756
rect 159416 11716 205088 11744
rect 159416 11704 159422 11716
rect 205082 11704 205088 11716
rect 205140 11704 205146 11756
rect 267734 11704 267740 11756
rect 267792 11744 267798 11756
rect 488810 11744 488816 11756
rect 267792 11716 488816 11744
rect 267792 11704 267798 11716
rect 488810 11704 488816 11716
rect 488868 11704 488874 11756
rect 157978 10344 157984 10396
rect 158036 10384 158042 10396
rect 201586 10384 201592 10396
rect 158036 10356 201592 10384
rect 158036 10344 158042 10356
rect 201586 10344 201592 10356
rect 201644 10344 201650 10396
rect 252554 10344 252560 10396
rect 252612 10384 252618 10396
rect 448514 10384 448520 10396
rect 252612 10356 448520 10384
rect 252612 10344 252618 10356
rect 448514 10344 448520 10356
rect 448572 10344 448578 10396
rect 173158 10276 173164 10328
rect 173216 10316 173222 10328
rect 240134 10316 240140 10328
rect 173216 10288 240140 10316
rect 173216 10276 173222 10288
rect 240134 10276 240140 10288
rect 240192 10276 240198 10328
rect 266354 10276 266360 10328
rect 266412 10316 266418 10328
rect 484762 10316 484768 10328
rect 266412 10288 484768 10316
rect 266412 10276 266418 10288
rect 484762 10276 484768 10288
rect 484820 10276 484826 10328
rect 263594 8916 263600 8968
rect 263652 8956 263658 8968
rect 478138 8956 478144 8968
rect 263652 8928 478144 8956
rect 263652 8916 263658 8928
rect 478138 8916 478144 8928
rect 478196 8916 478202 8968
rect 234614 8100 234620 8152
rect 234672 8140 234678 8152
rect 403618 8140 403624 8152
rect 234672 8112 403624 8140
rect 234672 8100 234678 8112
rect 403618 8100 403624 8112
rect 403676 8100 403682 8152
rect 237374 8032 237380 8084
rect 237432 8072 237438 8084
rect 410794 8072 410800 8084
rect 237432 8044 410800 8072
rect 237432 8032 237438 8044
rect 410794 8032 410800 8044
rect 410852 8032 410858 8084
rect 242894 7964 242900 8016
rect 242952 8004 242958 8016
rect 424962 8004 424968 8016
rect 242952 7976 424968 8004
rect 242952 7964 242958 7976
rect 424962 7964 424968 7976
rect 425020 7964 425026 8016
rect 248414 7896 248420 7948
rect 248472 7936 248478 7948
rect 439130 7936 439136 7948
rect 248472 7908 439136 7936
rect 248472 7896 248478 7908
rect 439130 7896 439136 7908
rect 439188 7896 439194 7948
rect 251174 7828 251180 7880
rect 251232 7868 251238 7880
rect 446214 7868 446220 7880
rect 251232 7840 446220 7868
rect 251232 7828 251238 7840
rect 446214 7828 446220 7840
rect 446272 7828 446278 7880
rect 253934 7760 253940 7812
rect 253992 7800 253998 7812
rect 453298 7800 453304 7812
rect 253992 7772 453304 7800
rect 253992 7760 253998 7772
rect 453298 7760 453304 7772
rect 453356 7760 453362 7812
rect 256694 7692 256700 7744
rect 256752 7732 256758 7744
rect 460382 7732 460388 7744
rect 256752 7704 460388 7732
rect 256752 7692 256758 7704
rect 460382 7692 460388 7704
rect 460440 7692 460446 7744
rect 259454 7624 259460 7676
rect 259512 7664 259518 7676
rect 467466 7664 467472 7676
rect 259512 7636 467472 7664
rect 259512 7624 259518 7636
rect 467466 7624 467472 7636
rect 467524 7624 467530 7676
rect 156598 7556 156604 7608
rect 156656 7596 156662 7608
rect 197906 7596 197912 7608
rect 156656 7568 197912 7596
rect 156656 7556 156662 7568
rect 197906 7556 197912 7568
rect 197964 7556 197970 7608
rect 262214 7556 262220 7608
rect 262272 7596 262278 7608
rect 474550 7596 474556 7608
rect 262272 7568 474556 7596
rect 262272 7556 262278 7568
rect 474550 7556 474556 7568
rect 474608 7556 474614 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 120718 6848 120724 6860
rect 3476 6820 120724 6848
rect 3476 6808 3482 6820
rect 120718 6808 120724 6820
rect 120776 6808 120782 6860
rect 198734 6740 198740 6792
rect 198792 6780 198798 6792
rect 311434 6780 311440 6792
rect 198792 6752 311440 6780
rect 198792 6740 198798 6752
rect 311434 6740 311440 6752
rect 311492 6740 311498 6792
rect 200114 6672 200120 6724
rect 200172 6712 200178 6724
rect 315022 6712 315028 6724
rect 200172 6684 315028 6712
rect 200172 6672 200178 6684
rect 315022 6672 315028 6684
rect 315080 6672 315086 6724
rect 201494 6604 201500 6656
rect 201552 6644 201558 6656
rect 318518 6644 318524 6656
rect 201552 6616 318524 6644
rect 201552 6604 201558 6616
rect 318518 6604 318524 6616
rect 318576 6604 318582 6656
rect 202874 6536 202880 6588
rect 202932 6576 202938 6588
rect 322106 6576 322112 6588
rect 202932 6548 322112 6576
rect 202932 6536 202938 6548
rect 322106 6536 322112 6548
rect 322164 6536 322170 6588
rect 204254 6468 204260 6520
rect 204312 6508 204318 6520
rect 325602 6508 325608 6520
rect 204312 6480 325608 6508
rect 204312 6468 204318 6480
rect 325602 6468 325608 6480
rect 325660 6468 325666 6520
rect 205634 6400 205640 6452
rect 205692 6440 205698 6452
rect 329190 6440 329196 6452
rect 205692 6412 329196 6440
rect 205692 6400 205698 6412
rect 329190 6400 329196 6412
rect 329248 6400 329254 6452
rect 207014 6332 207020 6384
rect 207072 6372 207078 6384
rect 332686 6372 332692 6384
rect 207072 6344 332692 6372
rect 207072 6332 207078 6344
rect 332686 6332 332692 6344
rect 332744 6332 332750 6384
rect 208486 6264 208492 6316
rect 208544 6304 208550 6316
rect 336274 6304 336280 6316
rect 208544 6276 336280 6304
rect 208544 6264 208550 6276
rect 336274 6264 336280 6276
rect 336332 6264 336338 6316
rect 209774 6196 209780 6248
rect 209832 6236 209838 6248
rect 339862 6236 339868 6248
rect 209832 6208 339868 6236
rect 209832 6196 209838 6208
rect 339862 6196 339868 6208
rect 339920 6196 339926 6248
rect 142154 6128 142160 6180
rect 142212 6168 142218 6180
rect 166074 6168 166080 6180
rect 142212 6140 166080 6168
rect 142212 6128 142218 6140
rect 166074 6128 166080 6140
rect 166132 6128 166138 6180
rect 211246 6128 211252 6180
rect 211304 6168 211310 6180
rect 343358 6168 343364 6180
rect 211304 6140 343364 6168
rect 211304 6128 211310 6140
rect 343358 6128 343364 6140
rect 343416 6128 343422 6180
rect 173894 5380 173900 5432
rect 173952 5420 173958 5432
rect 247586 5420 247592 5432
rect 173952 5392 247592 5420
rect 173952 5380 173958 5392
rect 247586 5380 247592 5392
rect 247644 5380 247650 5432
rect 277394 5380 277400 5432
rect 277452 5420 277458 5432
rect 513558 5420 513564 5432
rect 277452 5392 513564 5420
rect 277452 5380 277458 5392
rect 513558 5380 513564 5392
rect 513616 5380 513622 5432
rect 175274 5312 175280 5364
rect 175332 5352 175338 5364
rect 251174 5352 251180 5364
rect 175332 5324 251180 5352
rect 175332 5312 175338 5324
rect 251174 5312 251180 5324
rect 251232 5312 251238 5364
rect 278774 5312 278780 5364
rect 278832 5352 278838 5364
rect 517146 5352 517152 5364
rect 278832 5324 517152 5352
rect 278832 5312 278838 5324
rect 517146 5312 517152 5324
rect 517204 5312 517210 5364
rect 176654 5244 176660 5296
rect 176712 5284 176718 5296
rect 254670 5284 254676 5296
rect 176712 5256 254676 5284
rect 176712 5244 176718 5256
rect 254670 5244 254676 5256
rect 254728 5244 254734 5296
rect 280154 5244 280160 5296
rect 280212 5284 280218 5296
rect 520734 5284 520740 5296
rect 280212 5256 520740 5284
rect 280212 5244 280218 5256
rect 520734 5244 520740 5256
rect 520792 5244 520798 5296
rect 178034 5176 178040 5228
rect 178092 5216 178098 5228
rect 258258 5216 258264 5228
rect 178092 5188 258264 5216
rect 178092 5176 178098 5188
rect 258258 5176 258264 5188
rect 258316 5176 258322 5228
rect 281534 5176 281540 5228
rect 281592 5216 281598 5228
rect 524230 5216 524236 5228
rect 281592 5188 524236 5216
rect 281592 5176 281598 5188
rect 524230 5176 524236 5188
rect 524288 5176 524294 5228
rect 179414 5108 179420 5160
rect 179472 5148 179478 5160
rect 261754 5148 261760 5160
rect 179472 5120 261760 5148
rect 179472 5108 179478 5120
rect 261754 5108 261760 5120
rect 261812 5108 261818 5160
rect 282914 5108 282920 5160
rect 282972 5148 282978 5160
rect 527818 5148 527824 5160
rect 282972 5120 527824 5148
rect 282972 5108 282978 5120
rect 527818 5108 527824 5120
rect 527876 5108 527882 5160
rect 180794 5040 180800 5092
rect 180852 5080 180858 5092
rect 265342 5080 265348 5092
rect 180852 5052 265348 5080
rect 180852 5040 180858 5052
rect 265342 5040 265348 5052
rect 265400 5040 265406 5092
rect 284294 5040 284300 5092
rect 284352 5080 284358 5092
rect 531314 5080 531320 5092
rect 284352 5052 531320 5080
rect 284352 5040 284358 5052
rect 531314 5040 531320 5052
rect 531372 5040 531378 5092
rect 182174 4972 182180 5024
rect 182232 5012 182238 5024
rect 268838 5012 268844 5024
rect 182232 4984 268844 5012
rect 182232 4972 182238 4984
rect 268838 4972 268844 4984
rect 268896 4972 268902 5024
rect 285674 4972 285680 5024
rect 285732 5012 285738 5024
rect 534902 5012 534908 5024
rect 285732 4984 534908 5012
rect 285732 4972 285738 4984
rect 534902 4972 534908 4984
rect 534960 4972 534966 5024
rect 183554 4904 183560 4956
rect 183612 4944 183618 4956
rect 272426 4944 272432 4956
rect 183612 4916 272432 4944
rect 183612 4904 183618 4916
rect 272426 4904 272432 4916
rect 272484 4904 272490 4956
rect 287054 4904 287060 4956
rect 287112 4944 287118 4956
rect 538398 4944 538404 4956
rect 287112 4916 538404 4944
rect 287112 4904 287118 4916
rect 538398 4904 538404 4916
rect 538456 4904 538462 4956
rect 184934 4836 184940 4888
rect 184992 4876 184998 4888
rect 276014 4876 276020 4888
rect 184992 4848 276020 4876
rect 184992 4836 184998 4848
rect 276014 4836 276020 4848
rect 276072 4836 276078 4888
rect 288434 4836 288440 4888
rect 288492 4876 288498 4888
rect 541986 4876 541992 4888
rect 288492 4848 541992 4876
rect 288492 4836 288498 4848
rect 541986 4836 541992 4848
rect 542044 4836 542050 4888
rect 140774 4768 140780 4820
rect 140832 4808 140838 4820
rect 162486 4808 162492 4820
rect 140832 4780 162492 4808
rect 140832 4768 140838 4780
rect 162486 4768 162492 4780
rect 162544 4768 162550 4820
rect 186314 4768 186320 4820
rect 186372 4808 186378 4820
rect 279510 4808 279516 4820
rect 186372 4780 279516 4808
rect 186372 4768 186378 4780
rect 279510 4768 279516 4780
rect 279568 4768 279574 4820
rect 289814 4768 289820 4820
rect 289872 4808 289878 4820
rect 545482 4808 545488 4820
rect 289872 4780 545488 4808
rect 289872 4768 289878 4780
rect 545482 4768 545488 4780
rect 545540 4768 545546 4820
rect 129826 4088 129832 4140
rect 129884 4128 129890 4140
rect 134150 4128 134156 4140
rect 129884 4100 134156 4128
rect 129884 4088 129890 4100
rect 134150 4088 134156 4100
rect 134208 4088 134214 4140
rect 136634 4088 136640 4140
rect 136692 4128 136698 4140
rect 151814 4128 151820 4140
rect 136692 4100 151820 4128
rect 136692 4088 136698 4100
rect 151814 4088 151820 4100
rect 151872 4088 151878 4140
rect 138014 4020 138020 4072
rect 138072 4060 138078 4072
rect 155402 4060 155408 4072
rect 138072 4032 155408 4060
rect 138072 4020 138078 4032
rect 155402 4020 155408 4032
rect 155460 4020 155466 4072
rect 139394 3952 139400 4004
rect 139452 3992 139458 4004
rect 158898 3992 158904 4004
rect 139452 3964 158904 3992
rect 139452 3952 139458 3964
rect 158898 3952 158904 3964
rect 158956 3952 158962 4004
rect 143534 3884 143540 3936
rect 143592 3924 143598 3936
rect 169570 3924 169576 3936
rect 143592 3896 169576 3924
rect 143592 3884 143598 3896
rect 169570 3884 169576 3896
rect 169628 3884 169634 3936
rect 144914 3816 144920 3868
rect 144972 3856 144978 3868
rect 173158 3856 173164 3868
rect 144972 3828 173164 3856
rect 144972 3816 144978 3828
rect 173158 3816 173164 3828
rect 173216 3816 173222 3868
rect 146294 3748 146300 3800
rect 146352 3788 146358 3800
rect 176654 3788 176660 3800
rect 146352 3760 176660 3788
rect 146352 3748 146358 3760
rect 176654 3748 176660 3760
rect 176712 3748 176718 3800
rect 203518 3748 203524 3800
rect 203576 3788 203582 3800
rect 286594 3788 286600 3800
rect 203576 3760 286600 3788
rect 203576 3748 203582 3760
rect 286594 3748 286600 3760
rect 286652 3748 286658 3800
rect 313918 3748 313924 3800
rect 313976 3788 313982 3800
rect 435542 3788 435548 3800
rect 313976 3760 435548 3788
rect 313976 3748 313982 3760
rect 435542 3748 435548 3760
rect 435600 3748 435606 3800
rect 147674 3680 147680 3732
rect 147732 3720 147738 3732
rect 180242 3720 180248 3732
rect 147732 3692 180248 3720
rect 147732 3680 147738 3692
rect 180242 3680 180248 3692
rect 180300 3680 180306 3732
rect 210418 3680 210424 3732
rect 210476 3720 210482 3732
rect 293678 3720 293684 3732
rect 210476 3692 293684 3720
rect 210476 3680 210482 3692
rect 293678 3680 293684 3692
rect 293736 3680 293742 3732
rect 320818 3680 320824 3732
rect 320876 3720 320882 3732
rect 456886 3720 456892 3732
rect 320876 3692 456892 3720
rect 320876 3680 320882 3692
rect 456886 3680 456892 3692
rect 456944 3680 456950 3732
rect 131114 3612 131120 3664
rect 131172 3652 131178 3664
rect 137646 3652 137652 3664
rect 131172 3624 137652 3652
rect 131172 3612 131178 3624
rect 137646 3612 137652 3624
rect 137704 3612 137710 3664
rect 149054 3612 149060 3664
rect 149112 3652 149118 3664
rect 183738 3652 183744 3664
rect 149112 3624 183744 3652
rect 149112 3612 149118 3624
rect 183738 3612 183744 3624
rect 183796 3612 183802 3664
rect 213178 3612 213184 3664
rect 213236 3652 213242 3664
rect 297266 3652 297272 3664
rect 213236 3624 297272 3652
rect 213236 3612 213242 3624
rect 297266 3612 297272 3624
rect 297324 3612 297330 3664
rect 323578 3612 323584 3664
rect 323636 3652 323642 3664
rect 471054 3652 471060 3664
rect 323636 3624 471060 3652
rect 323636 3612 323642 3624
rect 471054 3612 471060 3624
rect 471112 3612 471118 3664
rect 133966 3544 133972 3596
rect 134024 3584 134030 3596
rect 144730 3584 144736 3596
rect 134024 3556 144736 3584
rect 134024 3544 134030 3556
rect 144730 3544 144736 3556
rect 144788 3544 144794 3596
rect 150434 3544 150440 3596
rect 150492 3584 150498 3596
rect 187326 3584 187332 3596
rect 150492 3556 187332 3584
rect 150492 3544 150498 3556
rect 187326 3544 187332 3556
rect 187384 3544 187390 3596
rect 206278 3544 206284 3596
rect 206336 3584 206342 3596
rect 290182 3584 290188 3596
rect 206336 3556 290188 3584
rect 206336 3544 206342 3556
rect 290182 3544 290188 3556
rect 290240 3544 290246 3596
rect 330478 3544 330484 3596
rect 330536 3584 330542 3596
rect 582190 3584 582196 3596
rect 330536 3556 582196 3584
rect 330536 3544 330542 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 135312 3488 141372 3516
rect 135312 3476 135318 3488
rect 125686 3408 125692 3460
rect 125744 3448 125750 3460
rect 128170 3448 128176 3460
rect 125744 3420 128176 3448
rect 125744 3408 125750 3420
rect 128170 3408 128176 3420
rect 128228 3408 128234 3460
rect 132494 3408 132500 3460
rect 132552 3448 132558 3460
rect 141234 3448 141240 3460
rect 132552 3420 141240 3448
rect 132552 3408 132558 3420
rect 141234 3408 141240 3420
rect 141292 3408 141298 3460
rect 141344 3448 141372 3488
rect 151906 3476 151912 3528
rect 151964 3516 151970 3528
rect 190822 3516 190828 3528
rect 151964 3488 190828 3516
rect 151964 3476 151970 3488
rect 190822 3476 190828 3488
rect 190880 3476 190886 3528
rect 199378 3476 199384 3528
rect 199436 3516 199442 3528
rect 283098 3516 283104 3528
rect 199436 3488 283104 3516
rect 199436 3476 199442 3488
rect 283098 3476 283104 3488
rect 283156 3476 283162 3528
rect 331858 3476 331864 3528
rect 331916 3516 331922 3528
rect 583386 3516 583392 3528
rect 331916 3488 583392 3516
rect 331916 3476 331922 3488
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 148318 3448 148324 3460
rect 141344 3420 148324 3448
rect 148318 3408 148324 3420
rect 148376 3408 148382 3460
rect 153194 3408 153200 3460
rect 153252 3448 153258 3460
rect 194410 3448 194416 3460
rect 153252 3420 194416 3448
rect 153252 3408 153258 3420
rect 194410 3408 194416 3420
rect 194468 3408 194474 3460
rect 218054 3408 218060 3460
rect 218112 3448 218118 3460
rect 219250 3448 219256 3460
rect 218112 3420 219256 3448
rect 218112 3408 218118 3420
rect 219250 3408 219256 3420
rect 219308 3408 219314 3460
rect 300762 3448 300768 3460
rect 219406 3420 300768 3448
rect 214558 3340 214564 3392
rect 214616 3380 214622 3392
rect 219406 3380 219434 3420
rect 300762 3408 300768 3420
rect 300820 3408 300826 3460
rect 327718 3408 327724 3460
rect 327776 3448 327782 3460
rect 580994 3448 581000 3460
rect 327776 3420 581000 3448
rect 327776 3408 327782 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 214616 3352 219434 3380
rect 214616 3340 214622 3352
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 448514 3340 448520 3392
rect 448572 3380 448578 3392
rect 449802 3380 449808 3392
rect 448572 3352 449808 3380
rect 448572 3340 448578 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 349154 2320 349160 2372
rect 349212 2360 349218 2372
rect 350442 2360 350448 2372
rect 349212 2332 350448 2360
rect 349212 2320 349218 2332
rect 350442 2320 350448 2332
rect 350500 2320 350506 2372
rect 398834 2320 398840 2372
rect 398892 2360 398898 2372
rect 400122 2360 400128 2372
rect 398892 2332 400128 2360
rect 398892 2320 398898 2332
rect 400122 2320 400128 2332
rect 400180 2320 400186 2372
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 170312 700680 170364 700732
rect 178316 700680 178368 700732
rect 154120 700612 154172 700664
rect 178408 700612 178460 700664
rect 137836 700544 137888 700596
rect 178040 700544 178092 700596
rect 105452 700476 105504 700528
rect 178224 700476 178276 700528
rect 392584 700476 392636 700528
rect 429844 700476 429896 700528
rect 177396 700408 177448 700460
rect 283840 700408 283892 700460
rect 366364 700408 366416 700460
rect 413652 700408 413704 700460
rect 72976 700340 73028 700392
rect 178132 700340 178184 700392
rect 186964 700340 187016 700392
rect 218980 700340 219032 700392
rect 360844 700340 360896 700392
rect 462320 700340 462372 700392
rect 89168 700272 89220 700324
rect 176660 700272 176712 700324
rect 177304 700272 177356 700324
rect 348792 700272 348844 700324
rect 363604 700272 363656 700324
rect 478512 700272 478564 700324
rect 24308 699660 24360 699712
rect 26884 699660 26936 699712
rect 192484 696940 192536 696992
rect 580172 696940 580224 696992
rect 170864 685856 170916 685908
rect 192576 685856 192628 685908
rect 351000 685856 351052 685908
rect 378784 685856 378836 685908
rect 530952 685856 531004 685908
rect 536840 685856 536892 685908
rect 3424 683136 3476 683188
rect 18604 683136 18656 683188
rect 3516 670692 3568 670744
rect 18696 670692 18748 670744
rect 538864 670692 538916 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 31024 656888 31076 656940
rect 537484 643084 537536 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 3148 618264 3200 618316
rect 25504 618264 25556 618316
rect 538956 616836 539008 616888
rect 580172 616836 580224 616888
rect 192576 607860 192628 607912
rect 213920 607860 213972 607912
rect 378784 607860 378836 607912
rect 394700 607860 394752 607912
rect 213920 607316 213972 607368
rect 216680 607316 216732 607368
rect 394700 607180 394752 607232
rect 397184 607180 397236 607232
rect 3240 605820 3292 605872
rect 11704 605820 11756 605872
rect 66812 597456 66864 597508
rect 84200 597456 84252 597508
rect 397736 597456 397788 597508
rect 436008 597456 436060 597508
rect 74908 597388 74960 597440
rect 92480 597388 92532 597440
rect 399484 597388 399536 597440
rect 434628 597388 434680 597440
rect 68744 597320 68796 597372
rect 85580 597320 85632 597372
rect 397828 597320 397880 597372
rect 437112 597320 437164 597372
rect 66168 597252 66220 597304
rect 82820 597252 82872 597304
rect 395344 597252 395396 597304
rect 434720 597252 434772 597304
rect 39212 597184 39264 597236
rect 74908 597184 74960 597236
rect 77116 597184 77168 597236
rect 95240 597184 95292 597236
rect 256700 597184 256752 597236
rect 274640 597184 274692 597236
rect 426532 597184 426584 597236
rect 444380 597184 444432 597236
rect 68836 597116 68888 597168
rect 86960 597116 87012 597168
rect 214748 597116 214800 597168
rect 258080 597116 258132 597168
rect 276020 597116 276072 597168
rect 425612 597116 425664 597168
rect 443644 597116 443696 597168
rect 36912 597048 36964 597100
rect 78036 597048 78088 597100
rect 96620 597048 96672 597100
rect 139308 597048 139360 597100
rect 178960 597048 179012 597100
rect 243084 597048 243136 597100
rect 260840 597048 260892 597100
rect 424968 597048 425020 597100
rect 441988 597048 442040 597100
rect 39948 596980 40000 597032
rect 56600 596980 56652 597032
rect 69756 596980 69808 597032
rect 88340 596980 88392 597032
rect 126888 596980 126940 597032
rect 177948 596980 178000 597032
rect 219716 596980 219768 597032
rect 236000 596980 236052 597032
rect 244280 596980 244332 597032
rect 262220 596980 262272 597032
rect 399668 596980 399720 597032
rect 416780 596980 416832 597032
rect 434628 596980 434680 597032
rect 452660 596980 452712 597032
rect 39672 596912 39724 596964
rect 59360 596912 59412 596964
rect 70400 596912 70452 596964
rect 71320 596912 71372 596964
rect 89720 596912 89772 596964
rect 118608 596912 118660 596964
rect 178776 596912 178828 596964
rect 218888 596912 218940 596964
rect 236184 596912 236236 596964
rect 244372 596912 244424 596964
rect 245476 596912 245528 596964
rect 263692 596912 263744 596964
rect 399944 596912 399996 596964
rect 419540 596912 419592 596964
rect 436008 596912 436060 596964
rect 454040 596912 454092 596964
rect 39488 596844 39540 596896
rect 63224 596844 63276 596896
rect 81440 596844 81492 596896
rect 121368 596844 121420 596896
rect 182824 596844 182876 596896
rect 219072 596844 219124 596896
rect 237380 596844 237432 596896
rect 253940 596844 253992 596896
rect 254584 596844 254636 596896
rect 273260 596844 273312 596896
rect 326988 596844 327040 596896
rect 359004 596844 359056 596896
rect 398288 596844 398340 596896
rect 418160 596844 418212 596896
rect 437112 596844 437164 596896
rect 455420 596844 455472 596896
rect 39764 596776 39816 596828
rect 64236 596776 64288 596828
rect 82820 596776 82872 596828
rect 117228 596776 117280 596828
rect 178868 596776 178920 596828
rect 219256 596776 219308 596828
rect 238760 596776 238812 596828
rect 245660 596776 245712 596828
rect 246488 596776 246540 596828
rect 265072 596776 265124 596828
rect 324228 596776 324280 596828
rect 357900 596776 357952 596828
rect 398564 596776 398616 596828
rect 419540 596776 419592 596828
rect 38384 596708 38436 596760
rect 64880 596708 64932 596760
rect 66168 596708 66220 596760
rect 114468 596708 114520 596760
rect 178684 596708 178736 596760
rect 218980 596708 219032 596760
rect 240140 596708 240192 596760
rect 252100 596708 252152 596760
rect 270592 596708 270644 596760
rect 321468 596708 321520 596760
rect 359096 596708 359148 596760
rect 398104 596708 398156 596760
rect 420920 596708 420972 596760
rect 39396 596640 39448 596692
rect 66812 596640 66864 596692
rect 111708 596640 111760 596692
rect 177856 596640 177908 596692
rect 217968 596640 218020 596692
rect 241520 596640 241572 596692
rect 252192 596640 252244 596692
rect 269120 596640 269172 596692
rect 318708 596640 318760 596692
rect 357716 596640 357768 596692
rect 399760 596640 399812 596692
rect 423128 596776 423180 596828
rect 441620 596776 441672 596828
rect 39304 596572 39356 596624
rect 68836 596572 68888 596624
rect 124128 596572 124180 596624
rect 191104 596572 191156 596624
rect 219164 596572 219216 596624
rect 243084 596572 243136 596624
rect 248420 596572 248472 596624
rect 266360 596572 266412 596624
rect 314568 596572 314620 596624
rect 357532 596572 357584 596624
rect 398472 596572 398524 596624
rect 424968 596572 425020 596624
rect 428004 596572 428056 596624
rect 447232 596572 447284 596624
rect 37648 596504 37700 596556
rect 67640 596504 67692 596556
rect 68744 596504 68796 596556
rect 108948 596504 109000 596556
rect 180064 596504 180116 596556
rect 218796 596504 218848 596556
rect 244280 596504 244332 596556
rect 249892 596504 249944 596556
rect 267924 596504 267976 596556
rect 315948 596504 316000 596556
rect 359188 596504 359240 596556
rect 398380 596504 398432 596556
rect 425612 596504 425664 596556
rect 426440 596504 426492 596556
rect 427636 596504 427688 596556
rect 445852 596504 445904 596556
rect 37188 596436 37240 596488
rect 69756 596436 69808 596488
rect 76012 596436 76064 596488
rect 94044 596436 94096 596488
rect 106188 596436 106240 596488
rect 177764 596436 177816 596488
rect 214840 596436 214892 596488
rect 244372 596436 244424 596488
rect 247132 596436 247184 596488
rect 266360 596436 266412 596488
rect 311808 596436 311860 596488
rect 357624 596436 357676 596488
rect 399576 596436 399628 596488
rect 426532 596436 426584 596488
rect 429200 596436 429252 596488
rect 448520 596436 448572 596488
rect 37096 596368 37148 596420
rect 70400 596368 70452 596420
rect 71780 596368 71832 596420
rect 91100 596368 91152 596420
rect 102048 596368 102100 596420
rect 177580 596368 177632 596420
rect 215116 596368 215168 596420
rect 245660 596368 245712 596420
rect 253480 596368 253532 596420
rect 271880 596368 271932 596420
rect 309048 596368 309100 596420
rect 356612 596368 356664 596420
rect 431960 596368 432012 596420
rect 449992 596368 450044 596420
rect 73160 596300 73212 596352
rect 91192 596300 91244 596352
rect 99288 596300 99340 596352
rect 177672 596300 177724 596352
rect 219808 596300 219860 596352
rect 253940 596300 253992 596352
rect 306104 596300 306156 596352
rect 357440 596300 357492 596352
rect 433432 596300 433484 596352
rect 451280 596300 451332 596352
rect 37924 596232 37976 596284
rect 77116 596232 77168 596284
rect 96528 596232 96580 596284
rect 177488 596232 177540 596284
rect 215024 596232 215076 596284
rect 256700 596232 256752 596284
rect 303528 596232 303580 596284
rect 358912 596232 358964 596284
rect 430672 596232 430724 596284
rect 448520 596232 448572 596284
rect 39120 596164 39172 596216
rect 55404 596164 55456 596216
rect 91008 596164 91060 596216
rect 200764 596164 200816 596216
rect 255412 596164 255464 596216
rect 273260 596164 273312 596216
rect 296352 596164 296404 596216
rect 357808 596164 357860 596216
rect 399852 596164 399904 596216
rect 415400 596164 415452 596216
rect 437480 596164 437532 596216
rect 456800 596164 456852 596216
rect 216312 594736 216364 594788
rect 249892 594736 249944 594788
rect 390192 594736 390244 594788
rect 477500 594736 477552 594788
rect 218704 594668 218756 594720
rect 253480 594668 253532 594720
rect 389916 594668 389968 594720
rect 480260 594668 480312 594720
rect 217324 594600 217376 594652
rect 252100 594600 252152 594652
rect 387524 594600 387576 594652
rect 483020 594600 483072 594652
rect 214564 594532 214616 594584
rect 255412 594532 255464 594584
rect 387156 594532 387208 594584
rect 485780 594532 485832 594584
rect 214656 594464 214708 594516
rect 259460 594464 259512 594516
rect 387340 594464 387392 594516
rect 488540 594464 488592 594516
rect 214472 594396 214524 594448
rect 259552 594396 259604 594448
rect 387616 594396 387668 594448
rect 489920 594396 489972 594448
rect 219900 594328 219952 594380
rect 285680 594328 285732 594380
rect 387432 594328 387484 594380
rect 492680 594328 492732 594380
rect 212356 594260 212408 594312
rect 280160 594260 280212 594312
rect 387248 594260 387300 594312
rect 495440 594260 495492 594312
rect 36636 594192 36688 594244
rect 71780 594192 71832 594244
rect 210976 594192 211028 594244
rect 287060 594192 287112 594244
rect 387064 594192 387116 594244
rect 498200 594192 498252 594244
rect 35808 594124 35860 594176
rect 73160 594124 73212 594176
rect 215208 594124 215260 594176
rect 292580 594124 292632 594176
rect 387708 594124 387760 594176
rect 500960 594124 501012 594176
rect 36728 594056 36780 594108
rect 76012 594056 76064 594108
rect 212448 594056 212500 594108
rect 289820 594056 289872 594108
rect 386972 594056 387024 594108
rect 502340 594056 502392 594108
rect 214380 593988 214432 594040
rect 247132 593988 247184 594040
rect 390376 593988 390428 594040
rect 474740 593988 474792 594040
rect 216496 593920 216548 593972
rect 248420 593920 248472 593972
rect 390008 593920 390060 593972
rect 473360 593920 473412 593972
rect 219348 593852 219400 593904
rect 252192 593852 252244 593904
rect 395068 593852 395120 593904
rect 438860 593852 438912 593904
rect 398012 591948 398064 592000
rect 426440 591948 426492 592000
rect 399300 591880 399352 591932
rect 429200 591880 429252 591932
rect 397920 591812 397972 591864
rect 428004 591812 428056 591864
rect 398196 591744 398248 591796
rect 430672 591744 430724 591796
rect 399208 591676 399260 591728
rect 431960 591676 432012 591728
rect 399392 591608 399444 591660
rect 433432 591608 433484 591660
rect 395804 591540 395856 591592
rect 437480 591540 437532 591592
rect 395160 591472 395212 591524
rect 440332 591472 440384 591524
rect 384396 591404 384448 591456
rect 445760 591404 445812 591456
rect 384304 591336 384356 591388
rect 447140 591336 447192 591388
rect 384488 591268 384540 591320
rect 449900 591268 449952 591320
rect 188344 590656 188396 590708
rect 579620 590656 579672 590708
rect 38476 585760 38528 585812
rect 217140 585760 217192 585812
rect 37740 585148 37792 585200
rect 38476 585148 38528 585200
rect 2780 579912 2832 579964
rect 4896 579912 4948 579964
rect 193864 576852 193916 576904
rect 579620 576852 579672 576904
rect 170864 567128 170916 567180
rect 213920 567128 213972 567180
rect 351092 567128 351144 567180
rect 394700 567128 394752 567180
rect 3424 565836 3476 565888
rect 35164 565836 35216 565888
rect 530952 565836 531004 565888
rect 536840 565836 536892 565888
rect 142068 565700 142120 565752
rect 204076 565700 204128 565752
rect 136548 565632 136600 565684
rect 203892 565632 203944 565684
rect 133788 565564 133840 565616
rect 203800 565564 203852 565616
rect 131028 565496 131080 565548
rect 203708 565496 203760 565548
rect 88248 565428 88300 565480
rect 200948 565428 201000 565480
rect 86868 565360 86920 565412
rect 200856 565360 200908 565412
rect 84108 565292 84160 565344
rect 201040 565292 201092 565344
rect 81348 565224 81400 565276
rect 203984 565224 204036 565276
rect 78588 565156 78640 565208
rect 203616 565156 203668 565208
rect 77208 565088 77260 565140
rect 203524 565088 203576 565140
rect 214932 563728 214984 563780
rect 249800 563728 249852 563780
rect 37832 563660 37884 563712
rect 217232 563660 217284 563712
rect 39028 563252 39080 563304
rect 40040 563252 40092 563304
rect 537668 563048 537720 563100
rect 579896 563048 579948 563100
rect 3424 553392 3476 553444
rect 25596 553392 25648 553444
rect 544384 536800 544436 536852
rect 580172 536800 580224 536852
rect 3424 527824 3476 527876
rect 8944 527824 8996 527876
rect 541624 524424 541676 524476
rect 580172 524424 580224 524476
rect 537576 510620 537628 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 14464 500964 14516 501016
rect 374644 487772 374696 487824
rect 397184 487772 397236 487824
rect 39028 485256 39080 485308
rect 39672 485256 39724 485308
rect 39764 485256 39816 485308
rect 39764 485052 39816 485104
rect 38936 484916 38988 484968
rect 39948 484916 40000 484968
rect 540244 484372 540296 484424
rect 580172 484372 580224 484424
rect 38108 480020 38160 480072
rect 217600 480020 217652 480072
rect 38292 479952 38344 480004
rect 216864 479952 216916 480004
rect 38568 479884 38620 479936
rect 216680 479884 216732 479936
rect 38016 479816 38068 479868
rect 217140 479816 217192 479868
rect 37832 479748 37884 479800
rect 217416 479748 217468 479800
rect 216864 479476 216916 479528
rect 217508 479476 217560 479528
rect 216680 479340 216732 479392
rect 217784 479340 217836 479392
rect 39120 478864 39172 478916
rect 56048 478864 56100 478916
rect 218336 478932 218388 478984
rect 217232 478864 217284 478916
rect 217600 478864 217652 478916
rect 219716 478864 219768 478916
rect 236000 478864 236052 478916
rect 36636 478592 36688 478644
rect 72332 478592 72384 478644
rect 73804 478592 73856 478644
rect 39212 478524 39264 478576
rect 74632 478524 74684 478576
rect 77208 478524 77260 478576
rect 398380 478524 398432 478576
rect 425520 478524 425572 478576
rect 35808 478456 35860 478508
rect 73160 478456 73212 478508
rect 399576 478456 399628 478508
rect 426624 478456 426676 478508
rect 37924 478388 37976 478440
rect 76932 478388 76984 478440
rect 78588 478388 78640 478440
rect 398012 478388 398064 478440
rect 427820 478388 427872 478440
rect 36728 478320 36780 478372
rect 75828 478320 75880 478372
rect 78220 478320 78272 478372
rect 399300 478320 399352 478372
rect 430120 478320 430172 478372
rect 430580 478320 430632 478372
rect 36912 478252 36964 478304
rect 78128 478252 78180 478304
rect 397920 478252 397972 478304
rect 428556 478252 428608 478304
rect 430028 478252 430080 478304
rect 37004 478184 37056 478236
rect 79508 478184 79560 478236
rect 398196 478184 398248 478236
rect 431316 478184 431368 478236
rect 433248 478184 433300 478236
rect 36820 478116 36872 478168
rect 80612 478116 80664 478168
rect 82728 478116 82780 478168
rect 399208 478116 399260 478168
rect 432512 478116 432564 478168
rect 434628 478116 434680 478168
rect 394332 477912 394384 477964
rect 398380 477912 398432 477964
rect 394424 477844 394476 477896
rect 399576 477844 399628 477896
rect 397276 477776 397328 477828
rect 399300 477776 399352 477828
rect 394516 477708 394568 477760
rect 398012 477708 398064 477760
rect 398288 477708 398340 477760
rect 400128 477708 400180 477760
rect 394608 477640 394660 477692
rect 397920 477640 397972 477692
rect 398472 477640 398524 477692
rect 424140 477640 424192 477692
rect 426164 477640 426216 477692
rect 397184 477572 397236 477624
rect 398104 477572 398156 477624
rect 399024 477572 399076 477624
rect 399484 477572 399536 477624
rect 397368 477504 397420 477556
rect 398196 477504 398248 477556
rect 398748 477504 398800 477556
rect 399208 477504 399260 477556
rect 399392 477504 399444 477556
rect 434444 477504 434496 477556
rect 436008 477572 436060 477624
rect 37096 477436 37148 477488
rect 70860 477436 70912 477488
rect 86960 477436 87012 477488
rect 87604 477436 87656 477488
rect 216496 477436 216548 477488
rect 217048 477436 217100 477488
rect 217324 477436 217376 477488
rect 252376 477436 252428 477488
rect 252468 477436 252520 477488
rect 269120 477436 269172 477488
rect 433432 477436 433484 477488
rect 434536 477436 434588 477488
rect 37188 477368 37240 477420
rect 70216 477368 70268 477420
rect 85580 477368 85632 477420
rect 86316 477368 86368 477420
rect 214380 477368 214432 477420
rect 214564 477368 214616 477420
rect 255320 477368 255372 477420
rect 260840 477368 260892 477420
rect 278780 477368 278832 477420
rect 433248 477368 433300 477420
rect 448520 477368 448572 477420
rect 37648 477300 37700 477352
rect 67640 477300 67692 477352
rect 39304 477232 39356 477284
rect 68744 477232 68796 477284
rect 39396 477164 39448 477216
rect 66536 477164 66588 477216
rect 67548 477164 67600 477216
rect 38384 477096 38436 477148
rect 64880 477096 64932 477148
rect 78588 477300 78640 477352
rect 95792 477300 95844 477352
rect 96528 477300 96580 477352
rect 78128 477232 78180 477284
rect 96988 477232 97040 477284
rect 214748 477300 214800 477352
rect 215116 477300 215168 477352
rect 245936 477300 245988 477352
rect 247132 477300 247184 477352
rect 266360 477300 266412 477352
rect 436008 477300 436060 477352
rect 452660 477300 452712 477352
rect 214840 477232 214892 477284
rect 245476 477232 245528 477284
rect 263600 477232 263652 477284
rect 263692 477232 263744 477284
rect 277676 477232 277728 477284
rect 430028 477232 430080 477284
rect 447140 477232 447192 477284
rect 85580 477164 85632 477216
rect 207020 477164 207072 477216
rect 208308 477164 208360 477216
rect 217048 477164 217100 477216
rect 219348 477164 219400 477216
rect 251272 477164 251324 477216
rect 252468 477164 252520 477216
rect 259368 477164 259420 477216
rect 276020 477164 276072 477216
rect 399668 477164 399720 477216
rect 416780 477164 416832 477216
rect 430580 477164 430632 477216
rect 448520 477164 448572 477216
rect 39764 477028 39816 477080
rect 63500 477028 63552 477080
rect 77208 477096 77260 477148
rect 93032 477096 93084 477148
rect 216404 477096 216456 477148
rect 250076 477096 250128 477148
rect 251088 477096 251140 477148
rect 255320 477096 255372 477148
rect 273260 477096 273312 477148
rect 399852 477096 399904 477148
rect 415400 477096 415452 477148
rect 427728 477096 427780 477148
rect 445760 477096 445812 477148
rect 86960 477028 87012 477080
rect 96528 477028 96580 477080
rect 215024 477028 215076 477080
rect 256976 477028 257028 477080
rect 274640 477028 274692 477080
rect 399944 477028 399996 477080
rect 419540 477028 419592 477080
rect 426624 477028 426676 477080
rect 444380 477028 444432 477080
rect 445668 477028 445720 477080
rect 458180 477028 458232 477080
rect 39488 476960 39540 477012
rect 63224 476960 63276 477012
rect 39580 476892 39632 476944
rect 60740 476892 60792 476944
rect 39028 476824 39080 476876
rect 59452 476824 59504 476876
rect 70860 476960 70912 477012
rect 89720 476960 89772 477012
rect 217968 476960 218020 477012
rect 218796 476960 218848 477012
rect 244280 476960 244332 477012
rect 252376 476960 252428 477012
rect 270500 476960 270552 477012
rect 399484 476960 399536 477012
rect 400128 476960 400180 477012
rect 418160 476960 418212 477012
rect 435732 476960 435784 477012
rect 454040 476960 454092 477012
rect 70216 476892 70268 476944
rect 88708 476892 88760 476944
rect 81808 476824 81860 476876
rect 82636 476824 82688 476876
rect 91100 476892 91152 476944
rect 92204 476892 92256 476944
rect 245936 476892 245988 476944
rect 264980 476892 265032 476944
rect 326988 476892 327040 476944
rect 359648 476892 359700 476944
rect 398840 476892 398892 476944
rect 399576 476892 399628 476944
rect 419540 476892 419592 476944
rect 437480 476892 437532 476944
rect 438124 476892 438176 476944
rect 456800 476892 456852 476944
rect 216404 476824 216456 476876
rect 218704 476824 218756 476876
rect 219256 476824 219308 476876
rect 253388 476824 253440 476876
rect 271880 476824 271932 476876
rect 324228 476824 324280 476876
rect 356980 476824 357032 476876
rect 399760 476824 399812 476876
rect 39672 476756 39724 476808
rect 58164 476756 58216 476808
rect 63500 476756 63552 476808
rect 64236 476756 64288 476808
rect 82820 476756 82872 476808
rect 83924 476756 83976 476808
rect 89720 476756 89772 476808
rect 218060 476756 218112 476808
rect 219348 476756 219400 476808
rect 220728 476756 220780 476808
rect 254492 476756 254544 476808
rect 273260 476756 273312 476808
rect 321468 476756 321520 476808
rect 359372 476756 359424 476808
rect 397184 476756 397236 476808
rect 420920 476756 420972 476808
rect 436836 476824 436888 476876
rect 455420 476824 455472 476876
rect 423128 476756 423180 476808
rect 441620 476756 441672 476808
rect 444196 476756 444248 476808
rect 456892 476756 456944 476808
rect 39856 476688 39908 476740
rect 57888 476688 57940 476740
rect 64880 476688 64932 476740
rect 84016 476688 84068 476740
rect 211712 476688 211764 476740
rect 219164 476688 219216 476740
rect 243176 476688 243228 476740
rect 260840 476688 260892 476740
rect 318708 476688 318760 476740
rect 359556 476688 359608 476740
rect 425520 476688 425572 476740
rect 443000 476688 443052 476740
rect 67548 476620 67600 476672
rect 85304 476620 85356 476672
rect 91284 476620 91336 476672
rect 78220 476552 78272 476604
rect 73160 476484 73212 476536
rect 91100 476484 91152 476536
rect 73804 476416 73856 476468
rect 93032 476484 93084 476536
rect 219808 476484 219860 476536
rect 220728 476484 220780 476536
rect 94412 476416 94464 476468
rect 210608 476416 210660 476468
rect 214564 476416 214616 476468
rect 216496 476416 216548 476468
rect 217048 476416 217100 476468
rect 91192 476348 91244 476400
rect 207020 476348 207072 476400
rect 214380 476348 214432 476400
rect 84016 476280 84068 476332
rect 210792 476280 210844 476332
rect 214840 476280 214892 476332
rect 248604 476620 248656 476672
rect 266360 476620 266412 476672
rect 315948 476620 316000 476672
rect 358176 476620 358228 476672
rect 434444 476620 434496 476672
rect 451372 476620 451424 476672
rect 251088 476552 251140 476604
rect 268200 476552 268252 476604
rect 314568 476552 314620 476604
rect 359464 476552 359516 476604
rect 395804 476552 395856 476604
rect 437480 476552 437532 476604
rect 244280 476484 244332 476536
rect 262220 476484 262272 476536
rect 311808 476484 311860 476536
rect 358084 476484 358136 476536
rect 397828 476484 397880 476536
rect 436836 476484 436888 476536
rect 309048 476416 309100 476468
rect 357164 476416 357216 476468
rect 426164 476416 426216 476468
rect 441988 476416 442040 476468
rect 306104 476348 306156 476400
rect 360200 476348 360252 476400
rect 397736 476348 397788 476400
rect 435732 476348 435784 476400
rect 303528 476280 303580 476332
rect 360292 476280 360344 476332
rect 434628 476280 434680 476332
rect 449900 476280 449952 476332
rect 91192 476212 91244 476264
rect 91284 476212 91336 476264
rect 213460 476212 213512 476264
rect 215116 476212 215168 476264
rect 217784 476212 217836 476264
rect 247132 476212 247184 476264
rect 302148 476212 302200 476264
rect 361672 476212 361724 476264
rect 394056 476212 394108 476264
rect 397736 476212 397788 476264
rect 398932 476212 398984 476264
rect 399668 476212 399720 476264
rect 82636 476144 82688 476196
rect 211712 476144 211764 476196
rect 214748 476144 214800 476196
rect 216404 476144 216456 476196
rect 259368 476144 259420 476196
rect 299388 476144 299440 476196
rect 359280 476144 359332 476196
rect 394148 476144 394200 476196
rect 395804 476144 395856 476196
rect 399208 476144 399260 476196
rect 399852 476144 399904 476196
rect 83924 476076 83976 476128
rect 217968 476076 218020 476128
rect 296260 476076 296312 476128
rect 357992 476076 358044 476128
rect 394240 476076 394292 476128
rect 397828 476076 397880 476128
rect 399300 476076 399352 476128
rect 399760 476076 399812 476128
rect 400128 476076 400180 476128
rect 433340 476076 433392 476128
rect 3056 474716 3108 474768
rect 7564 474716 7616 474768
rect 215852 474648 215904 474700
rect 268016 474648 268068 474700
rect 393964 474648 394016 474700
rect 395068 474648 395120 474700
rect 395436 474648 395488 474700
rect 477500 474648 477552 474700
rect 219072 474580 219124 474632
rect 273260 474580 273312 474632
rect 395620 474580 395672 474632
rect 480536 474580 480588 474632
rect 215944 474512 215996 474564
rect 270500 474512 270552 474564
rect 395712 474512 395764 474564
rect 483020 474512 483072 474564
rect 219716 474444 219768 474496
rect 276020 474444 276072 474496
rect 395804 474444 395856 474496
rect 485780 474444 485832 474496
rect 214840 474376 214892 474428
rect 277584 474376 277636 474428
rect 395988 474376 396040 474428
rect 488540 474376 488592 474428
rect 219624 474308 219676 474360
rect 285680 474308 285732 474360
rect 395896 474308 395948 474360
rect 490472 474308 490524 474360
rect 213092 474240 213144 474292
rect 280160 474240 280212 474292
rect 395252 474240 395304 474292
rect 492680 474240 492732 474292
rect 215760 474172 215812 474224
rect 282920 474172 282972 474224
rect 399484 474172 399536 474224
rect 502340 474172 502392 474224
rect 218704 474104 218756 474156
rect 292580 474104 292632 474156
rect 392400 474104 392452 474156
rect 495440 474104 495492 474156
rect 208952 474036 209004 474088
rect 287704 474036 287756 474088
rect 393044 474036 393096 474088
rect 498200 474036 498252 474088
rect 210332 473968 210384 474020
rect 289820 473968 289872 474020
rect 392952 473968 393004 474020
rect 500960 473968 501012 474020
rect 216036 473900 216088 473952
rect 264980 473900 265032 473952
rect 395528 473900 395580 473952
rect 474740 473900 474792 473952
rect 216220 473832 216272 473884
rect 263600 473832 263652 473884
rect 397920 473832 397972 473884
rect 465080 473832 465132 473884
rect 216312 473764 216364 473816
rect 260840 473764 260892 473816
rect 395068 473764 395120 473816
rect 438860 473764 438912 473816
rect 395160 471928 395212 471980
rect 440240 471928 440292 471980
rect 392492 471452 392544 471504
rect 445760 471452 445812 471504
rect 393228 471384 393280 471436
rect 447140 471384 447192 471436
rect 392768 471316 392820 471368
rect 449900 471316 449952 471368
rect 393136 471248 393188 471300
rect 505100 471248 505152 471300
rect 393872 471180 393924 471232
rect 395160 471180 395212 471232
rect 182916 470568 182968 470620
rect 580172 470568 580224 470620
rect 3516 462340 3568 462392
rect 15844 462340 15896 462392
rect 188436 456764 188488 456816
rect 580172 456764 580224 456816
rect 358820 454724 358872 454776
rect 359740 454724 359792 454776
rect 538220 454724 538272 454776
rect 216772 454656 216824 454708
rect 217692 454656 217744 454708
rect 396448 454656 396500 454708
rect 396632 454656 396684 454708
rect 179052 453296 179104 453348
rect 358820 453296 358872 453348
rect 214564 451868 214616 451920
rect 249800 451868 249852 451920
rect 216956 450780 217008 450832
rect 217324 450780 217376 450832
rect 217324 450508 217376 450560
rect 396540 450508 396592 450560
rect 210148 449216 210200 449268
rect 247040 449216 247092 449268
rect 71688 449148 71740 449200
rect 212540 449148 212592 449200
rect 3148 448536 3200 448588
rect 14556 448536 14608 448588
rect 142068 448468 142120 448520
rect 209228 448468 209280 448520
rect 139308 448400 139360 448452
rect 209412 448400 209464 448452
rect 136548 448332 136600 448384
rect 209044 448332 209096 448384
rect 133788 448264 133840 448316
rect 209596 448264 209648 448316
rect 131028 448196 131080 448248
rect 209504 448196 209556 448248
rect 91008 448128 91060 448180
rect 206560 448128 206612 448180
rect 88248 448060 88300 448112
rect 206652 448060 206704 448112
rect 86868 447992 86920 448044
rect 206744 447992 206796 448044
rect 84108 447924 84160 447976
rect 206468 447924 206520 447976
rect 81348 447856 81400 447908
rect 206376 447856 206428 447908
rect 78588 447788 78640 447840
rect 206284 447788 206336 447840
rect 143448 447720 143500 447772
rect 209320 447720 209372 447772
rect 146208 447652 146260 447704
rect 209136 447652 209188 447704
rect 170864 447040 170916 447092
rect 180156 447040 180208 447092
rect 351092 447040 351144 447092
rect 374644 447040 374696 447092
rect 530492 446972 530544 447024
rect 536840 446972 536892 447024
rect 218980 446360 219032 446412
rect 252560 446360 252612 446412
rect 124128 445680 124180 445732
rect 212264 445680 212316 445732
rect 121368 445612 121420 445664
rect 212172 445612 212224 445664
rect 118608 445544 118660 445596
rect 211988 445544 212040 445596
rect 117228 445476 117280 445528
rect 211804 445476 211856 445528
rect 114468 445408 114520 445460
rect 211896 445408 211948 445460
rect 106188 445340 106240 445392
rect 215024 445340 215076 445392
rect 104808 445272 104860 445324
rect 214472 445272 214524 445324
rect 102048 445204 102100 445256
rect 214288 445204 214340 445256
rect 99288 445136 99340 445188
rect 214748 445136 214800 445188
rect 96528 445068 96580 445120
rect 214656 445068 214708 445120
rect 68928 445000 68980 445052
rect 208584 445000 208636 445052
rect 126888 444932 126940 444984
rect 212080 444932 212132 444984
rect 129648 444864 129700 444916
rect 209688 444864 209740 444916
rect 178500 444320 178552 444372
rect 179052 444320 179104 444372
rect 77208 443640 77260 443692
rect 219900 443640 219952 443692
rect 38476 443232 38528 443284
rect 178500 443232 178552 443284
rect 548524 430584 548576 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 10324 422288 10376 422340
rect 540336 404336 540388 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 11796 397468 11848 397520
rect 217600 393320 217652 393372
rect 218060 393320 218112 393372
rect 217324 392028 217376 392080
rect 218704 392028 218756 392080
rect 218520 391960 218572 392012
rect 218704 391892 218756 391944
rect 547144 378156 547196 378208
rect 580172 378156 580224 378208
rect 3332 371220 3384 371272
rect 10416 371220 10468 371272
rect 362224 367140 362276 367192
rect 396724 367140 396776 367192
rect 358268 367072 358320 367124
rect 396540 367072 396592 367124
rect 396448 367004 396500 367056
rect 396724 367004 396776 367056
rect 543004 364352 543056 364404
rect 579804 364352 579856 364404
rect 38200 360000 38252 360052
rect 218612 360000 218664 360052
rect 224224 360000 224276 360052
rect 234068 360000 234120 360052
rect 396632 360000 396684 360052
rect 218520 359932 218572 359984
rect 210976 359864 211028 359916
rect 270500 359864 270552 359916
rect 311716 359864 311768 359916
rect 357900 359864 357952 359916
rect 212448 359796 212500 359848
rect 273444 359796 273496 359848
rect 279332 359796 279384 359848
rect 357808 359796 357860 359848
rect 361580 359796 361632 359848
rect 362224 359796 362276 359848
rect 393780 359796 393832 359848
rect 394148 359796 394200 359848
rect 215208 359728 215260 359780
rect 276388 359728 276440 359780
rect 300676 359728 300728 359780
rect 395252 359728 395304 359780
rect 210332 359660 210384 359712
rect 273076 359660 273128 359712
rect 277124 359660 277176 359712
rect 398012 359660 398064 359712
rect 208952 359592 209004 359644
rect 270132 359592 270184 359644
rect 271236 359592 271288 359644
rect 397828 359592 397880 359644
rect 215760 359524 215812 359576
rect 263508 359524 263560 359576
rect 264612 359524 264664 359576
rect 398196 359524 398248 359576
rect 213092 359456 213144 359508
rect 259736 359456 259788 359508
rect 261300 359456 261352 359508
rect 398564 359456 398616 359508
rect 217324 359388 217376 359440
rect 276112 359388 276164 359440
rect 314292 359388 314344 359440
rect 359648 359388 359700 359440
rect 219624 359320 219676 359372
rect 266820 359320 266872 359372
rect 397368 359320 397420 359372
rect 211068 359252 211120 359304
rect 257252 359252 257304 359304
rect 214840 359184 214892 359236
rect 256884 359184 256936 359236
rect 397276 359116 397328 359168
rect 217232 358708 217284 358760
rect 396816 358708 396868 358760
rect 216956 358640 217008 358692
rect 217324 358640 217376 358692
rect 397092 358640 397144 358692
rect 217876 358572 217928 358624
rect 396908 358572 396960 358624
rect 218336 358504 218388 358556
rect 236000 358504 236052 358556
rect 305460 358504 305512 358556
rect 359556 358504 359608 358556
rect 216036 358436 216088 358488
rect 239956 358436 240008 358488
rect 302516 358436 302568 358488
rect 358176 358436 358228 358488
rect 215852 358368 215904 358420
rect 243636 358368 243688 358420
rect 302884 358368 302936 358420
rect 359188 358368 359240 358420
rect 215944 358300 215996 358352
rect 246948 358300 247000 358352
rect 299572 358300 299624 358352
rect 359464 358300 359516 358352
rect 147588 358232 147640 358284
rect 178408 358232 178460 358284
rect 219072 358232 219124 358284
rect 250260 358232 250312 358284
rect 296628 358232 296680 358284
rect 358084 358232 358136 358284
rect 146852 358164 146904 358216
rect 178316 358164 178368 358216
rect 219716 358164 219768 358216
rect 253572 358164 253624 358216
rect 293684 358164 293736 358216
rect 357164 358164 357216 358216
rect 146484 358096 146536 358148
rect 186964 358096 187016 358148
rect 216220 358096 216272 358148
rect 235908 358096 235960 358148
rect 236000 358096 236052 358148
rect 399208 358096 399260 358148
rect 38476 358028 38528 358080
rect 200120 358028 200172 358080
rect 216128 358028 216180 358080
rect 227812 358028 227864 358080
rect 216312 357960 216364 358012
rect 231860 357960 231912 358012
rect 218704 357892 218756 357944
rect 230020 357892 230072 357944
rect 397000 358028 397052 358080
rect 416044 358028 416096 358080
rect 308404 357960 308456 358012
rect 359372 357960 359424 358012
rect 311348 357892 311400 357944
rect 356980 357892 357032 357944
rect 218888 357824 218940 357876
rect 223396 357824 223448 357876
rect 314660 357824 314712 357876
rect 359004 357824 359056 357876
rect 3332 357416 3384 357468
rect 36544 357416 36596 357468
rect 262128 357348 262180 357400
rect 399300 357348 399352 357400
rect 423128 357348 423180 357400
rect 423588 357348 423640 357400
rect 262772 357280 262824 357332
rect 398196 357280 398248 357332
rect 398656 357280 398708 357332
rect 398840 357280 398892 357332
rect 399116 357280 399168 357332
rect 433432 357280 433484 357332
rect 263600 357212 263652 357264
rect 263968 357212 264020 357264
rect 394240 357212 394292 357264
rect 268292 357144 268344 357196
rect 268568 357144 268620 357196
rect 397368 357144 397420 357196
rect 399024 357144 399076 357196
rect 434628 357144 434680 357196
rect 444288 357212 444340 357264
rect 456800 357212 456852 357264
rect 451464 357144 451516 357196
rect 394056 357076 394108 357128
rect 394424 357076 394476 357128
rect 436008 357076 436060 357128
rect 445668 357076 445720 357128
rect 458180 357076 458232 357128
rect 266360 357008 266412 357060
rect 267556 357008 267608 357060
rect 394608 357008 394660 357060
rect 243544 356940 243596 356992
rect 262128 356940 262180 356992
rect 265072 356940 265124 356992
rect 265716 356940 265768 356992
rect 398380 357008 398432 357060
rect 398748 357008 398800 357060
rect 431960 357008 432012 357060
rect 449992 357008 450044 357060
rect 257344 356872 257396 356924
rect 275928 356872 275980 356924
rect 428556 356940 428608 356992
rect 436008 356940 436060 356992
rect 454040 356940 454092 356992
rect 394332 356872 394384 356924
rect 394608 356872 394660 356924
rect 397276 356872 397328 356924
rect 430672 356872 430724 356924
rect 434628 356872 434680 356924
rect 452752 356872 452804 356924
rect 491944 356872 491996 356924
rect 498200 356872 498252 356924
rect 251272 356804 251324 356856
rect 269764 356804 269816 356856
rect 270408 356804 270460 356856
rect 272156 356804 272208 356856
rect 398840 356804 398892 356856
rect 436836 356804 436888 356856
rect 455420 356804 455472 356856
rect 249708 356736 249760 356788
rect 266360 356736 266412 356788
rect 266452 356736 266504 356788
rect 394516 356736 394568 356788
rect 252100 356668 252152 356720
rect 254584 356668 254636 356720
rect 273352 356668 273404 356720
rect 274456 356668 274508 356720
rect 398196 356668 398248 356720
rect 424968 356668 425020 356720
rect 60648 356600 60700 356652
rect 62764 356600 62816 356652
rect 244924 356600 244976 356652
rect 262772 356600 262824 356652
rect 274548 356600 274600 356652
rect 394424 356600 394476 356652
rect 394608 356600 394660 356652
rect 426900 356600 426952 356652
rect 250076 356532 250128 356584
rect 268292 356532 268344 356584
rect 275928 356532 275980 356584
rect 394148 356532 394200 356584
rect 394240 356532 394292 356584
rect 425428 356532 425480 356584
rect 426348 356532 426400 356584
rect 437572 356736 437624 356788
rect 438400 356736 438452 356788
rect 456800 356736 456852 356788
rect 429200 356668 429252 356720
rect 430028 356668 430080 356720
rect 448520 356668 448572 356720
rect 428556 356600 428608 356652
rect 447140 356600 447192 356652
rect 464436 356600 464488 356652
rect 467840 356600 467892 356652
rect 427636 356532 427688 356584
rect 445760 356532 445812 356584
rect 258816 356464 258868 356516
rect 277032 356464 277084 356516
rect 393780 356464 393832 356516
rect 394608 356464 394660 356516
rect 423588 356464 423640 356516
rect 441712 356464 441764 356516
rect 471244 356464 471296 356516
rect 477500 356464 477552 356516
rect 255320 356396 255372 356448
rect 255780 356396 255832 356448
rect 274548 356396 274600 356448
rect 397368 356396 397420 356448
rect 429200 356396 429252 356448
rect 430672 356396 430724 356448
rect 448520 356396 448572 356448
rect 251456 356328 251508 356380
rect 252284 356328 252336 356380
rect 271144 356328 271196 356380
rect 398380 356328 398432 356380
rect 426348 356328 426400 356380
rect 443000 356328 443052 356380
rect 479524 356328 479576 356380
rect 488540 356328 488592 356380
rect 77208 356260 77260 356312
rect 196532 356260 196584 356312
rect 244280 356260 244332 356312
rect 245568 356260 245620 356312
rect 263600 356260 263652 356312
rect 270408 356260 270460 356312
rect 397276 356260 397328 356312
rect 426900 356260 426952 356312
rect 444380 356260 444432 356312
rect 467196 356260 467248 356312
rect 474740 356260 474792 356312
rect 476764 356260 476816 356312
rect 483020 356260 483072 356312
rect 494704 356260 494756 356312
rect 500960 356260 501012 356312
rect 68928 356192 68980 356244
rect 192116 356192 192168 356244
rect 245660 356192 245712 356244
rect 246856 356192 246908 356244
rect 265072 356192 265124 356244
rect 274456 356192 274508 356244
rect 399024 356192 399076 356244
rect 424968 356192 425020 356244
rect 441988 356192 442040 356244
rect 482284 356192 482336 356244
rect 489920 356192 489972 356244
rect 74080 356124 74132 356176
rect 203156 356124 203208 356176
rect 233700 356124 233752 356176
rect 248696 356124 248748 356176
rect 249708 356124 249760 356176
rect 252836 356124 252888 356176
rect 253388 356124 253440 356176
rect 272156 356124 272208 356176
rect 394148 356124 394200 356176
rect 436836 356124 436888 356176
rect 472716 356124 472768 356176
rect 480536 356124 480588 356176
rect 487804 356124 487856 356176
rect 495440 356124 495492 356176
rect 64328 356056 64380 356108
rect 65524 356056 65576 356108
rect 68928 356056 68980 356108
rect 198372 356056 198424 356108
rect 247132 356056 247184 356108
rect 266452 356056 266504 356108
rect 394608 356056 394660 356108
rect 437572 356056 437624 356108
rect 457444 356056 457496 356108
rect 460940 356056 460992 356108
rect 467104 356056 467156 356108
rect 470784 356056 470836 356108
rect 476856 356056 476908 356108
rect 492680 356056 492732 356108
rect 497464 356056 497516 356108
rect 505100 356056 505152 356108
rect 210516 355988 210568 356040
rect 260196 355988 260248 356040
rect 210700 355920 210752 355972
rect 260104 355920 260156 355972
rect 210608 355852 210660 355904
rect 255320 355852 255372 355904
rect 208308 355784 208360 355836
rect 251456 355784 251508 355836
rect 216404 355716 216456 355768
rect 258816 355716 258868 355768
rect 215116 355648 215168 355700
rect 257344 355648 257396 355700
rect 210792 355580 210844 355632
rect 244280 355580 244332 355632
rect 275652 355580 275704 355632
rect 292580 355580 292632 355632
rect 310980 355580 311032 355632
rect 322940 355580 322992 355632
rect 217600 355512 217652 355564
rect 251272 355512 251324 355564
rect 290740 355512 290792 355564
rect 360200 355512 360252 355564
rect 216496 355444 216548 355496
rect 250076 355444 250128 355496
rect 287796 355444 287848 355496
rect 360292 355444 360344 355496
rect 219256 355376 219308 355428
rect 251088 355376 251140 355428
rect 284852 355376 284904 355428
rect 361672 355376 361724 355428
rect 39028 355308 39080 355360
rect 199844 355308 199896 355360
rect 217784 355308 217836 355360
rect 247132 355308 247184 355360
rect 281908 355308 281960 355360
rect 359280 355308 359332 355360
rect 218796 355240 218848 355292
rect 238116 355240 238168 355292
rect 239588 355240 239640 355292
rect 264980 355240 265032 355292
rect 217416 355172 217468 355224
rect 230388 355172 230440 355224
rect 210424 355104 210476 355156
rect 225236 355104 225288 355156
rect 251088 354696 251140 354748
rect 252836 354696 252888 354748
rect 278964 354628 279016 354680
rect 357992 354628 358044 354680
rect 309508 354560 309560 354612
rect 392952 354560 393004 354612
rect 306564 354492 306616 354544
rect 393044 354492 393096 354544
rect 303620 354424 303672 354476
rect 392400 354424 392452 354476
rect 297732 354356 297784 354408
rect 395896 354356 395948 354408
rect 294788 354288 294840 354340
rect 395988 354288 396040 354340
rect 291844 354220 291896 354272
rect 395804 354220 395856 354272
rect 269764 354152 269816 354204
rect 287060 354152 287112 354204
rect 288900 354152 288952 354204
rect 395712 354152 395764 354204
rect 285956 354084 286008 354136
rect 395620 354084 395672 354136
rect 283012 354016 283064 354068
rect 395436 354016 395488 354068
rect 38844 353948 38896 354000
rect 198740 353948 198792 354000
rect 218428 353948 218480 354000
rect 226340 353948 226392 354000
rect 231492 353948 231544 354000
rect 260840 353948 260892 354000
rect 280068 353948 280120 354000
rect 395528 353948 395580 354000
rect 288164 353880 288216 353932
rect 358912 353880 358964 353932
rect 291108 353812 291160 353864
rect 357440 353812 357492 353864
rect 313924 353744 313976 353796
rect 325700 353744 325752 353796
rect 219808 353200 219860 353252
rect 252100 353200 252152 353252
rect 38936 352520 38988 352572
rect 197636 352520 197688 352572
rect 215760 352520 215812 352572
rect 238760 352520 238812 352572
rect 191196 351908 191248 351960
rect 580172 351908 580224 351960
rect 213368 351840 213420 351892
rect 237012 351840 237064 351892
rect 280436 351840 280488 351892
rect 390376 351840 390428 351892
rect 210884 351772 210936 351824
rect 215760 351772 215812 351824
rect 216404 351772 216456 351824
rect 253204 351772 253256 351824
rect 276020 351772 276072 351824
rect 277492 351772 277544 351824
rect 390008 351772 390060 351824
rect 274548 351704 274600 351756
rect 389732 351704 389784 351756
rect 271604 351636 271656 351688
rect 390284 351636 390336 351688
rect 268292 351568 268344 351620
rect 390468 351568 390520 351620
rect 264980 351500 265032 351552
rect 390100 351500 390152 351552
rect 261668 351432 261720 351484
rect 389824 351432 389876 351484
rect 251732 351364 251784 351416
rect 392860 351364 392912 351416
rect 225328 351296 225380 351348
rect 245660 351296 245712 351348
rect 248052 351296 248104 351348
rect 392768 351296 392820 351348
rect 244740 351228 244792 351280
rect 393228 351228 393280 351280
rect 38384 351160 38436 351212
rect 191380 351160 191432 351212
rect 241060 351160 241112 351212
rect 392492 351160 392544 351212
rect 283380 351092 283432 351144
rect 390192 351092 390244 351144
rect 312452 351024 312504 351076
rect 399484 351024 399536 351076
rect 315396 350956 315448 351008
rect 393136 350956 393188 351008
rect 212724 350548 212776 350600
rect 213368 350548 213420 350600
rect 213460 350480 213512 350532
rect 225328 350480 225380 350532
rect 225604 350480 225656 350532
rect 248788 350480 248840 350532
rect 251088 350480 251140 350532
rect 93400 349800 93452 349852
rect 202972 349800 203024 349852
rect 247684 349800 247736 349852
rect 449900 349800 449952 349852
rect 217048 349052 217100 349104
rect 233700 349052 233752 349104
rect 303988 349052 304040 349104
rect 387248 349052 387300 349104
rect 301044 348984 301096 349036
rect 387432 348984 387484 349036
rect 298100 348916 298152 348968
rect 387616 348916 387668 348968
rect 295156 348848 295208 348900
rect 387340 348848 387392 348900
rect 292212 348780 292264 348832
rect 387156 348780 387208 348832
rect 289268 348712 289320 348764
rect 387524 348712 387576 348764
rect 286324 348644 286376 348696
rect 389916 348644 389968 348696
rect 248420 348576 248472 348628
rect 384488 348576 384540 348628
rect 76012 348508 76064 348560
rect 205364 348508 205416 348560
rect 245108 348508 245160 348560
rect 384304 348508 384356 348560
rect 14556 348440 14608 348492
rect 154948 348440 155000 348492
rect 241428 348440 241480 348492
rect 384396 348440 384448 348492
rect 134340 348372 134392 348424
rect 580448 348372 580500 348424
rect 306932 348304 306984 348356
rect 387064 348304 387116 348356
rect 309876 348236 309928 348288
rect 387708 348236 387760 348288
rect 312820 348168 312872 348220
rect 386972 348168 387024 348220
rect 78496 347080 78548 347132
rect 206100 347080 206152 347132
rect 133604 347012 133656 347064
rect 540336 347012 540388 347064
rect 140228 345652 140280 345704
rect 558920 345652 558972 345704
rect 3332 345040 3384 345092
rect 148324 345040 148376 345092
rect 212356 344972 212408 345024
rect 243544 344972 243596 345024
rect 211712 344564 211764 344616
rect 212356 344564 212408 344616
rect 73068 344360 73120 344412
rect 202420 344360 202472 344412
rect 244372 344360 244424 344412
rect 447232 344360 447284 344412
rect 136916 344292 136968 344344
rect 537668 344292 537720 344344
rect 257344 342932 257396 342984
rect 258264 342932 258316 342984
rect 38568 342864 38620 342916
rect 207940 342864 207992 342916
rect 228548 342864 228600 342916
rect 437480 342864 437532 342916
rect 213184 342184 213236 342236
rect 238024 342184 238076 342236
rect 81256 341640 81308 341692
rect 207572 341640 207624 341692
rect 237748 341640 237800 341692
rect 250076 341640 250128 341692
rect 18696 341572 18748 341624
rect 150900 341572 150952 341624
rect 236644 341572 236696 341624
rect 443092 341572 443144 341624
rect 142436 341504 142488 341556
rect 392584 341504 392636 341556
rect 211160 340892 211212 340944
rect 213184 340892 213236 340944
rect 216772 340824 216824 340876
rect 217968 340824 218020 340876
rect 244924 340824 244976 340876
rect 36544 340280 36596 340332
rect 157616 340280 157668 340332
rect 77024 340212 77076 340264
rect 204628 340212 204680 340264
rect 227444 340212 227496 340264
rect 258172 340212 258224 340264
rect 139124 340144 139176 340196
rect 538864 340144 538916 340196
rect 139860 338716 139912 338768
rect 580264 338716 580316 338768
rect 224868 337424 224920 337476
rect 395344 337424 395396 337476
rect 61384 337356 61436 337408
rect 195428 337356 195480 337408
rect 250996 337356 251048 337408
rect 452660 337356 452712 337408
rect 7564 335996 7616 336048
rect 154580 335996 154632 336048
rect 240692 335996 240744 336048
rect 445852 335996 445904 336048
rect 4896 333276 4948 333328
rect 152372 333276 152424 333328
rect 141700 333208 141752 333260
rect 360844 333208 360896 333260
rect 4804 331848 4856 331900
rect 151268 331848 151320 331900
rect 224132 331848 224184 331900
rect 434720 331848 434772 331900
rect 63408 330624 63460 330676
rect 192852 330624 192904 330676
rect 223028 330624 223080 330676
rect 255412 330624 255464 330676
rect 3516 330556 3568 330608
rect 156420 330556 156472 330608
rect 215300 330556 215352 330608
rect 430580 330556 430632 330608
rect 143540 330488 143592 330540
rect 364340 330488 364392 330540
rect 70308 329128 70360 329180
rect 200580 329128 200632 329180
rect 284484 329128 284536 329180
rect 300860 329128 300912 329180
rect 14464 329060 14516 329112
rect 153844 329060 153896 329112
rect 210884 329060 210936 329112
rect 427820 329060 427872 329112
rect 68836 327836 68888 327888
rect 199476 327836 199528 327888
rect 214196 327836 214248 327888
rect 249984 327836 250036 327888
rect 11796 327768 11848 327820
rect 156052 327768 156104 327820
rect 232596 327768 232648 327820
rect 440240 327768 440292 327820
rect 133236 327700 133288 327752
rect 543004 327700 543056 327752
rect 59268 326408 59320 326460
rect 192024 326408 192076 326460
rect 138020 326340 138072 326392
rect 538956 326340 539008 326392
rect 143172 324912 143224 324964
rect 366364 324912 366416 324964
rect 131764 324300 131816 324352
rect 580172 324300 580224 324352
rect 137652 323688 137704 323740
rect 193864 323688 193916 323740
rect 25596 323620 25648 323672
rect 152740 323620 152792 323672
rect 66168 323552 66220 323604
rect 195796 323552 195848 323604
rect 65524 322260 65576 322312
rect 194324 322260 194376 322312
rect 138388 322192 138440 322244
rect 537484 322192 537536 322244
rect 79968 320900 80020 320952
rect 206836 320900 206888 320952
rect 257620 320900 257672 320952
rect 457536 320900 457588 320952
rect 135076 320832 135128 320884
rect 540244 320832 540296 320884
rect 306196 319472 306248 319524
rect 491944 319472 491996 319524
rect 142068 319404 142120 319456
rect 363604 319404 363656 319456
rect 3332 318792 3384 318844
rect 87604 318792 87656 318844
rect 139492 318180 139544 318232
rect 192484 318180 192536 318232
rect 75828 318112 75880 318164
rect 203064 318112 203116 318164
rect 10324 318044 10376 318096
rect 155684 318044 155736 318096
rect 270868 318044 270920 318096
rect 464436 318044 464488 318096
rect 62028 316684 62080 316736
rect 196900 316684 196952 316736
rect 267556 316684 267608 316736
rect 464344 316684 464396 316736
rect 245476 315392 245528 315444
rect 251456 315392 251508 315444
rect 91008 315324 91060 315376
rect 202788 315324 202840 315376
rect 209780 315324 209832 315376
rect 247224 315324 247276 315376
rect 259828 315324 259880 315376
rect 280160 315324 280212 315376
rect 285588 315324 285640 315376
rect 472716 315324 472768 315376
rect 136548 315256 136600 315308
rect 541624 315256 541676 315308
rect 88248 313964 88300 314016
rect 202052 313964 202104 314016
rect 6920 313896 6972 313948
rect 149428 313896 149480 313948
rect 309140 313896 309192 313948
rect 494704 313896 494756 313948
rect 62764 312536 62816 312588
rect 193956 312536 194008 312588
rect 224500 312536 224552 312588
rect 370504 312536 370556 312588
rect 132132 311856 132184 311908
rect 580172 311856 580224 311908
rect 78588 311176 78640 311228
rect 198004 311176 198056 311228
rect 31024 311108 31076 311160
rect 150532 311108 150584 311160
rect 300308 311108 300360 311160
rect 476856 311108 476908 311160
rect 81348 309816 81400 309868
rect 199108 309816 199160 309868
rect 15844 309748 15896 309800
rect 155316 309748 155368 309800
rect 303252 309748 303304 309800
rect 487804 309748 487856 309800
rect 35164 308456 35216 308508
rect 153108 308456 153160 308508
rect 74356 308388 74408 308440
rect 195060 308388 195112 308440
rect 279700 308388 279752 308440
rect 467196 308388 467248 308440
rect 106188 307096 106240 307148
rect 207204 307096 207256 307148
rect 8944 307028 8996 307080
rect 153476 307028 153528 307080
rect 243268 307028 243320 307080
rect 267740 307028 267792 307080
rect 282644 307028 282696 307080
rect 471244 307028 471296 307080
rect 137284 305600 137336 305652
rect 188344 305600 188396 305652
rect 254308 305600 254360 305652
rect 454684 305600 454736 305652
rect 3424 304988 3476 305040
rect 90364 304988 90416 305040
rect 256516 304376 256568 304428
rect 277400 304376 277452 304428
rect 235540 304308 235592 304360
rect 263692 304308 263744 304360
rect 278596 304308 278648 304360
rect 295340 304308 295392 304360
rect 104808 304240 104860 304292
rect 206008 304240 206060 304292
rect 260932 304240 260984 304292
rect 457444 304240 457496 304292
rect 102048 302948 102100 303000
rect 205732 302948 205784 303000
rect 11704 302880 11756 302932
rect 151636 302880 151688 302932
rect 288532 302880 288584 302932
rect 476764 302880 476816 302932
rect 99288 301520 99340 301572
rect 204996 301520 205048 301572
rect 26884 301452 26936 301504
rect 149796 301452 149848 301504
rect 276756 301452 276808 301504
rect 472624 301452 472676 301504
rect 96528 300092 96580 300144
rect 204260 300092 204312 300144
rect 273812 300092 273864 300144
rect 467104 300092 467156 300144
rect 258724 299412 258776 299464
rect 262036 299412 262088 299464
rect 71596 298800 71648 298852
rect 193588 298800 193640 298852
rect 25504 298732 25556 298784
rect 152004 298732 152056 298784
rect 258356 298732 258408 298784
rect 356796 298732 356848 298784
rect 131396 298120 131448 298172
rect 580172 298120 580224 298172
rect 260196 298052 260248 298104
rect 265348 298052 265400 298104
rect 305092 297712 305144 297764
rect 317420 297712 317472 297764
rect 254676 297644 254728 297696
rect 356704 297644 356756 297696
rect 232964 297576 233016 297628
rect 357072 297576 357124 297628
rect 228916 297508 228968 297560
rect 356888 297508 356940 297560
rect 263140 297440 263192 297492
rect 282920 297440 282972 297492
rect 294420 297440 294472 297492
rect 479524 297440 479576 297492
rect 38752 297372 38804 297424
rect 196164 297372 196216 297424
rect 219716 297372 219768 297424
rect 433340 297372 433392 297424
rect 177948 296216 178000 296268
rect 290004 296216 290056 296268
rect 178960 296148 179012 296200
rect 304724 296148 304776 296200
rect 71688 296080 71740 296132
rect 201868 296080 201920 296132
rect 281540 296080 281592 296132
rect 298192 296080 298244 296132
rect 299204 296080 299256 296132
rect 313280 296080 313332 296132
rect 177212 296012 177264 296064
rect 310612 296012 310664 296064
rect 38660 295944 38712 295996
rect 194692 295944 194744 295996
rect 249892 295944 249944 295996
rect 273352 295944 273404 295996
rect 297364 295944 297416 295996
rect 482284 295944 482336 295996
rect 177856 295060 177908 295112
rect 272340 295060 272392 295112
rect 191104 294992 191156 295044
rect 287060 294992 287112 295044
rect 178684 294924 178736 294976
rect 275284 294924 275336 294976
rect 178868 294856 178920 294908
rect 278228 294856 278280 294908
rect 182824 294788 182876 294840
rect 284116 294788 284168 294840
rect 178776 294720 178828 294772
rect 281172 294720 281224 294772
rect 67548 294652 67600 294704
rect 197268 294652 197320 294704
rect 58624 294584 58676 294636
rect 193220 294584 193272 294636
rect 296260 294584 296312 294636
rect 310520 294584 310572 294636
rect 315028 294584 315080 294636
rect 497464 294584 497516 294636
rect 203984 293904 204036 293956
rect 231124 293904 231176 293956
rect 201040 293836 201092 293888
rect 235172 293836 235224 293888
rect 218612 293768 218664 293820
rect 252652 293768 252704 293820
rect 200856 293700 200908 293752
rect 239220 293700 239272 293752
rect 200948 293632 201000 293684
rect 242900 293632 242952 293684
rect 177764 293564 177816 293616
rect 266084 293564 266136 293616
rect 272708 293564 272760 293616
rect 289912 293564 289964 293616
rect 290372 293564 290424 293616
rect 305000 293564 305052 293616
rect 203708 293496 203760 293548
rect 295892 293496 295944 293548
rect 203800 293428 203852 293480
rect 298836 293428 298888 293480
rect 203892 293360 203944 293412
rect 301780 293360 301832 293412
rect 86868 293292 86920 293344
rect 201316 293292 201368 293344
rect 204076 293292 204128 293344
rect 307668 293292 307720 293344
rect 308036 293292 308088 293344
rect 320180 293292 320232 293344
rect 200764 293224 200816 293276
rect 246212 293224 246264 293276
rect 264244 293224 264296 293276
rect 462320 293224 462372 293276
rect 3424 292544 3476 292596
rect 89720 292544 89772 292596
rect 135444 292068 135496 292120
rect 182916 292068 182968 292120
rect 302148 292068 302200 292120
rect 314752 292068 314804 292120
rect 177580 292000 177632 292052
rect 259460 292000 259512 292052
rect 266452 292000 266504 292052
rect 285680 292000 285732 292052
rect 293316 292000 293368 292052
rect 307760 292000 307812 292052
rect 180064 291932 180116 291984
rect 269396 291932 269448 291984
rect 287428 291932 287480 291984
rect 302240 291932 302292 291984
rect 84108 291864 84160 291916
rect 200212 291864 200264 291916
rect 217508 291864 217560 291916
rect 358268 291864 358320 291916
rect 56508 291796 56560 291848
rect 191748 291796 191800 291848
rect 208308 291796 208360 291848
rect 236092 291796 236144 291848
rect 246580 291796 246632 291848
rect 270592 291796 270644 291848
rect 291476 291796 291528 291848
rect 485780 291796 485832 291848
rect 212172 291116 212224 291168
rect 283748 291116 283800 291168
rect 212264 291048 212316 291100
rect 286692 291048 286744 291100
rect 212080 290980 212132 291032
rect 289636 290980 289688 291032
rect 209688 290912 209740 290964
rect 292580 290912 292632 290964
rect 209504 290844 209556 290896
rect 295524 290844 295576 290896
rect 209596 290776 209648 290828
rect 298468 290776 298520 290828
rect 209044 290708 209096 290760
rect 301412 290708 301464 290760
rect 209412 290640 209464 290692
rect 304356 290640 304408 290692
rect 209228 290572 209280 290624
rect 307300 290572 307352 290624
rect 209320 290504 209372 290556
rect 310244 290504 310296 290556
rect 89720 290436 89772 290488
rect 158260 290436 158312 290488
rect 312084 290436 312136 290488
rect 502340 290436 502392 290488
rect 206560 290368 206612 290420
rect 245844 290368 245896 290420
rect 206652 290300 206704 290352
rect 242532 290300 242584 290352
rect 206744 290232 206796 290284
rect 238852 290232 238904 290284
rect 209136 290164 209188 290216
rect 313188 290164 313240 290216
rect 316684 289756 316736 289808
rect 396724 289756 396776 289808
rect 90364 289212 90416 289264
rect 158628 289212 158680 289264
rect 217324 289212 217376 289264
rect 225972 289212 226024 289264
rect 3516 289144 3568 289196
rect 154212 289144 154264 289196
rect 217692 289144 217744 289196
rect 242164 289144 242216 289196
rect 132868 289076 132920 289128
rect 547144 289076 547196 289128
rect 316132 289008 316184 289060
rect 316684 289008 316736 289060
rect 217876 288396 217928 288448
rect 221556 288396 221608 288448
rect 220820 287920 220872 287972
rect 240232 287920 240284 287972
rect 148324 287852 148376 287904
rect 157156 287852 157208 287904
rect 206468 287852 206520 287904
rect 234804 287852 234856 287904
rect 241796 287852 241848 287904
rect 251272 287852 251324 287904
rect 132592 287784 132644 287836
rect 191196 287784 191248 287836
rect 211896 287784 211948 287836
rect 274916 287784 274968 287836
rect 87604 287716 87656 287768
rect 157892 287716 157944 287768
rect 211804 287716 211856 287768
rect 277860 287716 277912 287768
rect 10416 287648 10468 287700
rect 156788 287648 156840 287700
rect 211988 287648 212040 287700
rect 280804 287648 280856 287700
rect 176752 287580 176804 287632
rect 319536 287580 319588 287632
rect 172980 287512 173032 287564
rect 319720 287512 319772 287564
rect 167092 287444 167144 287496
rect 449900 287444 449952 287496
rect 172612 287376 172664 287428
rect 458180 287376 458232 287428
rect 182916 287308 182968 287360
rect 471980 287308 472032 287360
rect 184388 287240 184440 287292
rect 474740 287240 474792 287292
rect 187332 287172 187384 287224
rect 478880 287172 478932 287224
rect 189540 287104 189592 287156
rect 484400 287104 484452 287156
rect 190644 287036 190696 287088
rect 485780 287036 485832 287088
rect 146116 286492 146168 286544
rect 201500 286492 201552 286544
rect 221464 286492 221516 286544
rect 244280 286492 244332 286544
rect 166908 286424 166960 286476
rect 364340 286424 364392 286476
rect 168840 286356 168892 286408
rect 368480 286356 368532 286408
rect 170680 286288 170732 286340
rect 374000 286288 374052 286340
rect 172428 286220 172480 286272
rect 378140 286220 378192 286272
rect 174360 286152 174412 286204
rect 383660 286152 383712 286204
rect 176200 286084 176252 286136
rect 387800 286084 387852 286136
rect 181352 286016 181404 286068
rect 402980 286016 403032 286068
rect 182456 285948 182508 286000
rect 404360 285948 404412 286000
rect 182824 285880 182876 285932
rect 407120 285880 407172 285932
rect 184296 285812 184348 285864
rect 412640 285812 412692 285864
rect 185768 285744 185820 285796
rect 416780 285744 416832 285796
rect 187240 285676 187292 285728
rect 422300 285676 422352 285728
rect 145656 285268 145708 285320
rect 177396 285268 177448 285320
rect 144552 285200 144604 285252
rect 177304 285200 177356 285252
rect 203524 285200 203576 285252
rect 222476 285200 222528 285252
rect 229928 285200 229980 285252
rect 247132 285200 247184 285252
rect 134984 285132 135036 285184
rect 188436 285132 188488 285184
rect 206376 285132 206428 285184
rect 230572 285132 230624 285184
rect 260104 285132 260156 285184
rect 268476 285132 268528 285184
rect 170312 285064 170364 285116
rect 371240 285064 371292 285116
rect 40040 284996 40092 285048
rect 149060 284996 149112 285048
rect 172152 284996 172204 285048
rect 376760 284996 376812 285048
rect 18604 284928 18656 284980
rect 149980 284928 150032 284980
rect 175832 284928 175884 284980
rect 386420 284928 386472 284980
rect 179236 284860 179288 284912
rect 396080 284860 396132 284912
rect 179880 284792 179932 284844
rect 397460 284792 397512 284844
rect 185400 284724 185452 284776
rect 414020 284724 414072 284776
rect 186872 284656 186924 284708
rect 419540 284656 419592 284708
rect 188344 284588 188396 284640
rect 423680 284588 423732 284640
rect 189448 284520 189500 284572
rect 426440 284520 426492 284572
rect 190276 284452 190328 284504
rect 429200 284452 429252 284504
rect 169668 284384 169720 284436
rect 436100 284384 436152 284436
rect 179144 284316 179196 284368
rect 448520 284316 448572 284368
rect 130568 283772 130620 283824
rect 321100 283772 321152 283824
rect 178316 283704 178368 283756
rect 380900 283704 380952 283756
rect 187792 283636 187844 283688
rect 393320 283636 393372 283688
rect 136088 283568 136140 283620
rect 537576 283568 537628 283620
rect 169760 283500 169812 283552
rect 433340 283500 433392 283552
rect 116676 283432 116728 283484
rect 161020 283432 161072 283484
rect 174912 283432 174964 283484
rect 580540 283432 580592 283484
rect 119528 283364 119580 283416
rect 160100 283364 160152 283416
rect 173808 283364 173860 283416
rect 580724 283364 580776 283416
rect 126152 283296 126204 283348
rect 538956 283296 539008 283348
rect 127256 283228 127308 283280
rect 540244 283228 540296 283280
rect 125416 283160 125468 283212
rect 538864 283160 538916 283212
rect 128268 283092 128320 283144
rect 543096 283092 543148 283144
rect 129464 283024 129516 283076
rect 544384 283024 544436 283076
rect 126520 282956 126572 283008
rect 543004 282956 543056 283008
rect 143448 282888 143500 282940
rect 580356 282888 580408 282940
rect 192024 282820 192076 282872
rect 192300 282820 192352 282872
rect 200120 282820 200172 282872
rect 200764 282820 200816 282872
rect 202972 282820 203024 282872
rect 203340 282820 203392 282872
rect 206008 282820 206060 282872
rect 206284 282820 206336 282872
rect 208584 282820 208636 282872
rect 208860 282820 208912 282872
rect 212540 282820 212592 282872
rect 213276 282820 213328 282872
rect 219900 282820 219952 282872
rect 222200 282820 222252 282872
rect 258264 282820 258316 282872
rect 258540 282820 258592 282872
rect 259736 282820 259788 282872
rect 260012 282820 260064 282872
rect 266636 282820 266688 282872
rect 267004 282820 267056 282872
rect 203064 282752 203116 282804
rect 203708 282752 203760 282804
rect 166264 282548 166316 282600
rect 178040 282548 178092 282600
rect 90364 282480 90416 282532
rect 162860 282480 162912 282532
rect 173716 282480 173768 282532
rect 178316 282480 178368 282532
rect 148968 282412 149020 282464
rect 176660 282412 176712 282464
rect 177948 282412 178000 282464
rect 187792 282412 187844 282464
rect 148232 282344 148284 282396
rect 178224 282344 178276 282396
rect 180248 282344 180300 282396
rect 187884 282344 187936 282396
rect 206376 282344 206428 282396
rect 226524 282344 226576 282396
rect 127624 282276 127676 282328
rect 143448 282276 143500 282328
rect 147496 282276 147548 282328
rect 178132 282276 178184 282328
rect 186136 282276 186188 282328
rect 191656 282276 191708 282328
rect 214656 282276 214708 282328
rect 252284 282276 252336 282328
rect 130200 282208 130252 282260
rect 173808 282208 173860 282260
rect 181720 282208 181772 282260
rect 319904 282208 319956 282260
rect 129096 282140 129148 282192
rect 174912 282140 174964 282192
rect 178408 282140 178460 282192
rect 320088 282140 320140 282192
rect 15844 282072 15896 282124
rect 165068 282072 165120 282124
rect 175004 282072 175056 282124
rect 318156 282072 318208 282124
rect 133788 282004 133840 282056
rect 163964 282004 164016 282056
rect 169576 282004 169628 282056
rect 314844 282004 314896 282056
rect 120908 281936 120960 281988
rect 158904 281936 158956 281988
rect 171416 281936 171468 281988
rect 319444 281936 319496 281988
rect 119620 281868 119672 281920
rect 119436 281800 119488 281852
rect 156236 281800 156288 281852
rect 158812 281868 158864 281920
rect 164332 281868 164384 281920
rect 170956 281868 171008 281920
rect 320916 281868 320968 281920
rect 159180 281800 159232 281852
rect 169208 281800 169260 281852
rect 321008 281800 321060 281852
rect 120816 281732 120868 281784
rect 162124 281732 162176 281784
rect 174728 281732 174780 281784
rect 459560 281732 459612 281784
rect 120724 281664 120776 281716
rect 164700 281664 164752 281716
rect 167736 281664 167788 281716
rect 453304 281664 453356 281716
rect 121276 281596 121328 281648
rect 124588 281596 124640 281648
rect 156236 281596 156288 281648
rect 160284 281596 160336 281648
rect 168104 281596 168156 281648
rect 169760 281596 169812 281648
rect 176568 281596 176620 281648
rect 462320 281596 462372 281648
rect 143448 281528 143500 281580
rect 160652 281528 160704 281580
rect 166632 281528 166684 281580
rect 179420 281528 179472 281580
rect 188712 281528 188764 281580
rect 481640 281528 481692 281580
rect 184756 281052 184808 281104
rect 318064 281052 318116 281104
rect 130936 280984 130988 281036
rect 318248 280984 318300 281036
rect 3516 280916 3568 280968
rect 133788 280916 133840 280968
rect 178040 280916 178092 280968
rect 431960 280916 432012 280968
rect 3792 280848 3844 280900
rect 143448 280848 143500 280900
rect 191656 280848 191708 280900
rect 476120 280848 476172 280900
rect 3700 280780 3752 280832
rect 162492 280780 162544 280832
rect 175096 280780 175148 280832
rect 185492 280780 185544 280832
rect 185584 280780 185636 280832
rect 580632 280780 580684 280832
rect 131028 280712 131080 280764
rect 321192 280712 321244 280764
rect 129556 280644 129608 280696
rect 319996 280644 320048 280696
rect 168196 280576 168248 280628
rect 367100 280576 367152 280628
rect 180708 280508 180760 280560
rect 400220 280508 400272 280560
rect 115296 280440 115348 280492
rect 159548 280440 159600 280492
rect 173624 280440 173676 280492
rect 440240 280440 440292 280492
rect 119344 280372 119396 280424
rect 163596 280372 163648 280424
rect 171784 280372 171836 280424
rect 438860 280372 438912 280424
rect 116584 280304 116636 280356
rect 161572 280304 161624 280356
rect 177304 280304 177356 280356
rect 115204 280236 115256 280288
rect 161756 280236 161808 280288
rect 185492 280304 185544 280356
rect 443000 280304 443052 280356
rect 445760 280236 445812 280288
rect 3608 280168 3660 280220
rect 163458 280168 163510 280220
rect 165666 280168 165718 280220
rect 511264 280168 511316 280220
rect 121368 280100 121420 280152
rect 124220 280100 124272 280152
rect 314844 279828 314896 279880
rect 491300 279828 491352 279880
rect 179420 279760 179472 279812
rect 361672 279760 361724 279812
rect 187884 279692 187936 279744
rect 467840 279692 467892 279744
rect 177672 279624 177724 279676
rect 390560 279624 390612 279676
rect 3424 279488 3476 279540
rect 158812 279556 158864 279608
rect 180616 279556 180668 279608
rect 183928 279556 183980 279608
rect 409880 279556 409932 279608
rect 505100 279488 505152 279540
rect 3332 267656 3384 267708
rect 120908 267656 120960 267708
rect 321192 259360 321244 259412
rect 579804 259360 579856 259412
rect 2964 255212 3016 255264
rect 115296 255212 115348 255264
rect 321100 245556 321152 245608
rect 580172 245556 580224 245608
rect 3332 241408 3384 241460
rect 119620 241408 119672 241460
rect 320088 233928 320140 233980
rect 465448 233928 465500 233980
rect 319444 233860 319496 233912
rect 494152 233860 494204 233912
rect 319996 233180 320048 233232
rect 579988 233180 580040 233232
rect 321008 232976 321060 233028
rect 453212 232976 453264 233028
rect 453304 232976 453356 233028
rect 489368 232976 489420 233028
rect 491944 232976 491996 233028
rect 503720 232976 503772 233028
rect 320916 232908 320968 232960
rect 455880 232908 455932 232960
rect 456064 232908 456116 232960
rect 520464 232908 520516 232960
rect 319904 232840 319956 232892
rect 469772 232840 469824 232892
rect 469864 232840 469916 232892
rect 525248 232840 525300 232892
rect 319720 232772 319772 232824
rect 496544 232772 496596 232824
rect 319536 232704 319588 232756
rect 501328 232704 501380 232756
rect 320824 232636 320876 232688
rect 508504 232636 508556 232688
rect 319812 232568 319864 232620
rect 510896 232568 510948 232620
rect 511264 232568 511316 232620
rect 527640 232568 527692 232620
rect 319628 232500 319680 232552
rect 522856 232500 522908 232552
rect 319444 231820 319496 231872
rect 537208 231820 537260 231872
rect 319536 230460 319588 230512
rect 530032 230460 530084 230512
rect 3056 215228 3108 215280
rect 119528 215228 119580 215280
rect 544384 206932 544436 206984
rect 580172 206932 580224 206984
rect 3332 188980 3384 189032
rect 119436 188980 119488 189032
rect 543096 166948 543148 167000
rect 580172 166948 580224 167000
rect 3056 164160 3108 164212
rect 116676 164160 116728 164212
rect 3332 150356 3384 150408
rect 115204 150356 115256 150408
rect 540336 139340 540388 139392
rect 579804 139340 579856 139392
rect 3332 137912 3384 137964
rect 116584 137912 116636 137964
rect 540244 126896 540296 126948
rect 580172 126896 580224 126948
rect 543004 113092 543056 113144
rect 579620 113092 579672 113144
rect 3332 111732 3384 111784
rect 120816 111732 120868 111784
rect 3332 97928 3384 97980
rect 90364 97928 90416 97980
rect 538956 86912 539008 86964
rect 580172 86912 580224 86964
rect 314108 80588 314160 80640
rect 318064 80588 318116 80640
rect 318248 78684 318300 78736
rect 358820 78684 358872 78736
rect 225788 78616 225840 78668
rect 231124 78616 231176 78668
rect 234068 78616 234120 78668
rect 239404 78616 239456 78668
rect 312728 78616 312780 78668
rect 318340 78616 318392 78668
rect 188528 78548 188580 78600
rect 199384 78548 199436 78600
rect 189908 78480 189960 78532
rect 203524 78480 203576 78532
rect 315488 78480 315540 78532
rect 319444 78480 319496 78532
rect 191288 78412 191340 78464
rect 206284 78412 206336 78464
rect 311348 78412 311400 78464
rect 319536 78412 319588 78464
rect 192668 78344 192720 78396
rect 210424 78344 210476 78396
rect 195428 78276 195480 78328
rect 214564 78276 214616 78328
rect 304448 78276 304500 78328
rect 327724 78276 327776 78328
rect 194048 78208 194100 78260
rect 213184 78208 213236 78260
rect 307208 78208 307260 78260
rect 331864 78208 331916 78260
rect 159548 78140 159600 78192
rect 208400 78140 208452 78192
rect 305828 78140 305880 78192
rect 330484 78140 330536 78192
rect 160928 78072 160980 78124
rect 211160 78072 211212 78124
rect 261668 78072 261720 78124
rect 323584 78072 323636 78124
rect 1400 78004 1452 78056
rect 123024 78004 123076 78056
rect 162308 78004 162360 78056
rect 215300 78004 215352 78056
rect 236828 78004 236880 78056
rect 242164 78004 242216 78056
rect 256148 78004 256200 78056
rect 320824 78004 320876 78056
rect 20 77936 72 77988
rect 121644 77936 121696 77988
rect 163688 77936 163740 77988
rect 218060 77936 218112 77988
rect 218888 77936 218940 77988
rect 228364 77936 228416 77988
rect 247868 77936 247920 77988
rect 313924 77936 313976 77988
rect 239588 77392 239640 77444
rect 244924 77392 244976 77444
rect 242348 77324 242400 77376
rect 246304 77324 246356 77376
rect 125048 77256 125100 77308
rect 125600 77256 125652 77308
rect 129188 77256 129240 77308
rect 129740 77256 129792 77308
rect 155408 77256 155460 77308
rect 156604 77256 156656 77308
rect 156788 77256 156840 77308
rect 157984 77256 158036 77308
rect 158168 77256 158220 77308
rect 159364 77256 159416 77308
rect 171968 77256 172020 77308
rect 173164 77256 173216 77308
rect 214748 77256 214800 77308
rect 217324 77256 217376 77308
rect 221648 77256 221700 77308
rect 224224 77256 224276 77308
rect 240968 77256 241020 77308
rect 242256 77256 242308 77308
rect 245108 77256 245160 77308
rect 247684 77256 247736 77308
rect 165068 75148 165120 75200
rect 222200 75148 222252 75200
rect 195980 73788 196032 73840
rect 303620 73788 303672 73840
rect 538956 73108 539008 73160
rect 579988 73108 580040 73160
rect 224224 48968 224276 49020
rect 367100 48968 367152 49020
rect 309140 48220 309192 48272
rect 494888 48220 494940 48272
rect 307760 48152 307812 48204
rect 361580 48152 361632 48204
rect 404912 48152 404964 48204
rect 121276 46860 121328 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 119344 45500 119396 45552
rect 212540 44888 212592 44940
rect 346400 44888 346452 44940
rect 242256 44820 242308 44872
rect 416780 44820 416832 44872
rect 227720 43460 227772 43512
rect 385040 43460 385092 43512
rect 168380 43392 168432 43444
rect 233240 43392 233292 43444
rect 300860 43392 300912 43444
rect 572720 43392 572772 43444
rect 271880 42032 271932 42084
rect 498200 42032 498252 42084
rect 264980 40672 265032 40724
rect 481640 40672 481692 40724
rect 231860 39380 231912 39432
rect 396080 39380 396132 39432
rect 296720 39312 296772 39364
rect 563060 39312 563112 39364
rect 222292 37952 222344 38004
rect 371240 37952 371292 38004
rect 245660 37884 245712 37936
rect 431960 37884 432012 37936
rect 215392 36524 215444 36576
rect 353300 36524 353352 36576
rect 216680 35164 216732 35216
rect 357440 35164 357492 35216
rect 230480 33736 230532 33788
rect 391940 33736 391992 33788
rect 229100 31016 229152 31068
rect 389180 31016 389232 31068
rect 226340 29656 226392 29708
rect 382280 29656 382332 29708
rect 302240 29588 302292 29640
rect 576860 29588 576912 29640
rect 244924 28296 244976 28348
rect 414020 28296 414072 28348
rect 276020 28228 276072 28280
rect 509240 28228 509292 28280
rect 231124 26936 231176 26988
rect 378140 26936 378192 26988
rect 299480 26868 299532 26920
rect 569960 26868 570012 26920
rect 223580 25576 223632 25628
rect 374000 25576 374052 25628
rect 298100 25508 298152 25560
rect 565820 25508 565872 25560
rect 242164 24148 242216 24200
rect 407120 24148 407172 24200
rect 292580 24080 292632 24132
rect 552020 24080 552072 24132
rect 239404 22788 239456 22840
rect 398840 22788 398892 22840
rect 295340 22720 295392 22772
rect 558920 22720 558972 22772
rect 219440 21428 219492 21480
rect 364340 21428 364392 21480
rect 293960 21360 294012 21412
rect 556160 21360 556212 21412
rect 3424 20612 3476 20664
rect 15844 20612 15896 20664
rect 121368 20612 121420 20664
rect 579988 20612 580040 20664
rect 217324 19932 217376 19984
rect 349160 19932 349212 19984
rect 228364 18640 228416 18692
rect 360200 18640 360252 18692
rect 172520 18572 172572 18624
rect 242992 18572 243044 18624
rect 291200 18572 291252 18624
rect 547880 18572 547932 18624
rect 247684 17280 247736 17332
rect 427820 17280 427872 17332
rect 274640 17212 274692 17264
rect 506480 17212 506532 17264
rect 258080 15920 258132 15972
rect 463976 15920 464028 15972
rect 169760 15852 169812 15904
rect 236552 15852 236604 15904
rect 273260 15852 273312 15904
rect 502984 15852 503036 15904
rect 246304 14492 246356 14544
rect 420920 14492 420972 14544
rect 167000 14424 167052 14476
rect 229376 14424 229428 14476
rect 270500 14424 270552 14476
rect 495440 14424 495492 14476
rect 249800 13132 249852 13184
rect 442632 13132 442684 13184
rect 165620 13064 165672 13116
rect 226340 13064 226392 13116
rect 269120 13064 269172 13116
rect 492312 13064 492364 13116
rect 197360 11772 197412 11824
rect 307944 11772 307996 11824
rect 159364 11704 159416 11756
rect 205088 11704 205140 11756
rect 267740 11704 267792 11756
rect 488816 11704 488868 11756
rect 157984 10344 158036 10396
rect 201592 10344 201644 10396
rect 252560 10344 252612 10396
rect 448520 10344 448572 10396
rect 173164 10276 173216 10328
rect 240140 10276 240192 10328
rect 266360 10276 266412 10328
rect 484768 10276 484820 10328
rect 263600 8916 263652 8968
rect 478144 8916 478196 8968
rect 234620 8100 234672 8152
rect 403624 8100 403676 8152
rect 237380 8032 237432 8084
rect 410800 8032 410852 8084
rect 242900 7964 242952 8016
rect 424968 7964 425020 8016
rect 248420 7896 248472 7948
rect 439136 7896 439188 7948
rect 251180 7828 251232 7880
rect 446220 7828 446272 7880
rect 253940 7760 253992 7812
rect 453304 7760 453356 7812
rect 256700 7692 256752 7744
rect 460388 7692 460440 7744
rect 259460 7624 259512 7676
rect 467472 7624 467524 7676
rect 156604 7556 156656 7608
rect 197912 7556 197964 7608
rect 262220 7556 262272 7608
rect 474556 7556 474608 7608
rect 3424 6808 3476 6860
rect 120724 6808 120776 6860
rect 198740 6740 198792 6792
rect 311440 6740 311492 6792
rect 200120 6672 200172 6724
rect 315028 6672 315080 6724
rect 201500 6604 201552 6656
rect 318524 6604 318576 6656
rect 202880 6536 202932 6588
rect 322112 6536 322164 6588
rect 204260 6468 204312 6520
rect 325608 6468 325660 6520
rect 205640 6400 205692 6452
rect 329196 6400 329248 6452
rect 207020 6332 207072 6384
rect 332692 6332 332744 6384
rect 208492 6264 208544 6316
rect 336280 6264 336332 6316
rect 209780 6196 209832 6248
rect 339868 6196 339920 6248
rect 142160 6128 142212 6180
rect 166080 6128 166132 6180
rect 211252 6128 211304 6180
rect 343364 6128 343416 6180
rect 173900 5380 173952 5432
rect 247592 5380 247644 5432
rect 277400 5380 277452 5432
rect 513564 5380 513616 5432
rect 175280 5312 175332 5364
rect 251180 5312 251232 5364
rect 278780 5312 278832 5364
rect 517152 5312 517204 5364
rect 176660 5244 176712 5296
rect 254676 5244 254728 5296
rect 280160 5244 280212 5296
rect 520740 5244 520792 5296
rect 178040 5176 178092 5228
rect 258264 5176 258316 5228
rect 281540 5176 281592 5228
rect 524236 5176 524288 5228
rect 179420 5108 179472 5160
rect 261760 5108 261812 5160
rect 282920 5108 282972 5160
rect 527824 5108 527876 5160
rect 180800 5040 180852 5092
rect 265348 5040 265400 5092
rect 284300 5040 284352 5092
rect 531320 5040 531372 5092
rect 182180 4972 182232 5024
rect 268844 4972 268896 5024
rect 285680 4972 285732 5024
rect 534908 4972 534960 5024
rect 183560 4904 183612 4956
rect 272432 4904 272484 4956
rect 287060 4904 287112 4956
rect 538404 4904 538456 4956
rect 184940 4836 184992 4888
rect 276020 4836 276072 4888
rect 288440 4836 288492 4888
rect 541992 4836 542044 4888
rect 140780 4768 140832 4820
rect 162492 4768 162544 4820
rect 186320 4768 186372 4820
rect 279516 4768 279568 4820
rect 289820 4768 289872 4820
rect 545488 4768 545540 4820
rect 129832 4088 129884 4140
rect 134156 4088 134208 4140
rect 136640 4088 136692 4140
rect 151820 4088 151872 4140
rect 138020 4020 138072 4072
rect 155408 4020 155460 4072
rect 139400 3952 139452 4004
rect 158904 3952 158956 4004
rect 143540 3884 143592 3936
rect 169576 3884 169628 3936
rect 144920 3816 144972 3868
rect 173164 3816 173216 3868
rect 146300 3748 146352 3800
rect 176660 3748 176712 3800
rect 203524 3748 203576 3800
rect 286600 3748 286652 3800
rect 313924 3748 313976 3800
rect 435548 3748 435600 3800
rect 147680 3680 147732 3732
rect 180248 3680 180300 3732
rect 210424 3680 210476 3732
rect 293684 3680 293736 3732
rect 320824 3680 320876 3732
rect 456892 3680 456944 3732
rect 131120 3612 131172 3664
rect 137652 3612 137704 3664
rect 149060 3612 149112 3664
rect 183744 3612 183796 3664
rect 213184 3612 213236 3664
rect 297272 3612 297324 3664
rect 323584 3612 323636 3664
rect 471060 3612 471112 3664
rect 133972 3544 134024 3596
rect 144736 3544 144788 3596
rect 150440 3544 150492 3596
rect 187332 3544 187384 3596
rect 206284 3544 206336 3596
rect 290188 3544 290240 3596
rect 330484 3544 330536 3596
rect 582196 3544 582248 3596
rect 135260 3476 135312 3528
rect 125692 3408 125744 3460
rect 128176 3408 128228 3460
rect 132500 3408 132552 3460
rect 141240 3408 141292 3460
rect 151912 3476 151964 3528
rect 190828 3476 190880 3528
rect 199384 3476 199436 3528
rect 283104 3476 283156 3528
rect 331864 3476 331916 3528
rect 583392 3476 583444 3528
rect 148324 3408 148376 3460
rect 153200 3408 153252 3460
rect 194416 3408 194468 3460
rect 218060 3408 218112 3460
rect 219256 3408 219308 3460
rect 214564 3340 214616 3392
rect 300768 3408 300820 3460
rect 327724 3408 327776 3460
rect 581000 3408 581052 3460
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 448520 3340 448572 3392
rect 449808 3340 449860 3392
rect 349160 2320 349212 2372
rect 350448 2320 350500 2372
rect 398840 2320 398892 2372
rect 400128 2320 400180 2372
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 4804 632120 4856 632126
rect 2832 632088 2834 632097
rect 4804 632062 4856 632068
rect 2778 632023 2834 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 2778 580000 2834 580009
rect 2778 579935 2780 579944
rect 2832 579935 2834 579944
rect 2780 579906 2832 579912
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3424 527856
rect 3476 527847 3478 527856
rect 3424 527818 3476 527824
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3436 306374 3464 514791
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3514 410544 3570 410553
rect 3514 410479 3570 410488
rect 3528 330614 3556 410479
rect 4816 331906 4844 632062
rect 4896 579964 4948 579970
rect 4896 579906 4948 579912
rect 4908 333334 4936 579906
rect 4896 333328 4948 333334
rect 4896 333270 4948 333276
rect 4804 331900 4856 331906
rect 4804 331842 4856 331848
rect 3516 330608 3568 330614
rect 3516 330550 3568 330556
rect 6932 313954 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 699718 24348 703520
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 26884 699712 26936 699718
rect 26884 699654 26936 699660
rect 18604 683188 18656 683194
rect 18604 683130 18656 683136
rect 11704 605872 11756 605878
rect 11704 605814 11756 605820
rect 8944 527876 8996 527882
rect 8944 527818 8996 527824
rect 7564 474768 7616 474774
rect 7564 474710 7616 474716
rect 7576 336054 7604 474710
rect 7564 336048 7616 336054
rect 7564 335990 7616 335996
rect 6920 313948 6972 313954
rect 6920 313890 6972 313896
rect 8956 307086 8984 527818
rect 10324 422340 10376 422346
rect 10324 422282 10376 422288
rect 10336 318102 10364 422282
rect 10416 371272 10468 371278
rect 10416 371214 10468 371220
rect 10324 318096 10376 318102
rect 10324 318038 10376 318044
rect 8944 307080 8996 307086
rect 8944 307022 8996 307028
rect 3436 306346 3556 306374
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305046 3464 306167
rect 3424 305040 3476 305046
rect 3424 304982 3476 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3528 289202 3556 306346
rect 3516 289196 3568 289202
rect 3516 289138 3568 289144
rect 10428 287706 10456 371214
rect 11716 302938 11744 605814
rect 14464 501016 14516 501022
rect 14464 500958 14516 500964
rect 11796 397520 11848 397526
rect 11796 397462 11848 397468
rect 11808 327826 11836 397462
rect 14476 329118 14504 500958
rect 15844 462392 15896 462398
rect 15844 462334 15896 462340
rect 14556 448588 14608 448594
rect 14556 448530 14608 448536
rect 14568 348498 14596 448530
rect 14556 348492 14608 348498
rect 14556 348434 14608 348440
rect 14464 329112 14516 329118
rect 14464 329054 14516 329060
rect 11796 327820 11848 327826
rect 11796 327762 11848 327768
rect 15856 309806 15884 462334
rect 15844 309800 15896 309806
rect 15844 309742 15896 309748
rect 11704 302932 11756 302938
rect 11704 302874 11756 302880
rect 10416 287700 10468 287706
rect 10416 287642 10468 287648
rect 18616 284986 18644 683130
rect 18696 670744 18748 670750
rect 18696 670686 18748 670692
rect 18708 341630 18736 670686
rect 25504 618316 25556 618322
rect 25504 618258 25556 618264
rect 18696 341624 18748 341630
rect 18696 341566 18748 341572
rect 25516 298790 25544 618258
rect 25596 553444 25648 553450
rect 25596 553386 25648 553392
rect 25608 323678 25636 553386
rect 25596 323672 25648 323678
rect 25596 323614 25648 323620
rect 26896 301510 26924 699654
rect 40052 683346 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700398 73016 703520
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 89180 700330 89208 703520
rect 105464 700534 105492 703520
rect 137848 700602 137876 703520
rect 154132 700670 154160 703520
rect 170324 700738 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170312 700732 170364 700738
rect 170312 700674 170364 700680
rect 178316 700732 178368 700738
rect 178316 700674 178368 700680
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 137836 700596 137888 700602
rect 137836 700538 137888 700544
rect 178040 700596 178092 700602
rect 178040 700538 178092 700544
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 177396 700460 177448 700466
rect 177396 700402 177448 700408
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 176660 700324 176712 700330
rect 176660 700266 176712 700272
rect 177304 700324 177356 700330
rect 177304 700266 177356 700272
rect 170862 685944 170918 685953
rect 170862 685879 170864 685888
rect 170916 685879 170918 685888
rect 170864 685850 170916 685856
rect 39960 683318 40080 683346
rect 31024 656940 31076 656946
rect 31024 656882 31076 656888
rect 31036 311166 31064 656882
rect 37830 636304 37886 636313
rect 37830 636239 37886 636248
rect 36912 597100 36964 597106
rect 36912 597042 36964 597048
rect 36818 596864 36874 596873
rect 36818 596799 36874 596808
rect 36636 594244 36688 594250
rect 36636 594186 36688 594192
rect 35808 594176 35860 594182
rect 35808 594118 35860 594124
rect 35164 565888 35216 565894
rect 35164 565830 35216 565836
rect 31024 311160 31076 311166
rect 31024 311102 31076 311108
rect 35176 308514 35204 565830
rect 35820 478514 35848 594118
rect 36648 478650 36676 594186
rect 36728 594108 36780 594114
rect 36728 594050 36780 594056
rect 36636 478644 36688 478650
rect 36636 478586 36688 478592
rect 35808 478508 35860 478514
rect 35808 478450 35860 478456
rect 36740 478378 36768 594050
rect 36728 478372 36780 478378
rect 36728 478314 36780 478320
rect 36832 478174 36860 596799
rect 36924 478310 36952 597042
rect 37002 597000 37058 597009
rect 37002 596935 37058 596944
rect 36912 478304 36964 478310
rect 36912 478246 36964 478252
rect 37016 478242 37044 596935
rect 37648 596556 37700 596562
rect 37648 596498 37700 596504
rect 37188 596488 37240 596494
rect 37188 596430 37240 596436
rect 37096 596420 37148 596426
rect 37096 596362 37148 596368
rect 37004 478236 37056 478242
rect 37004 478178 37056 478184
rect 36820 478168 36872 478174
rect 36820 478110 36872 478116
rect 37108 477494 37136 596362
rect 37096 477488 37148 477494
rect 37096 477430 37148 477436
rect 37200 477426 37228 596430
rect 37188 477420 37240 477426
rect 37188 477362 37240 477368
rect 37660 477358 37688 596498
rect 37740 585200 37792 585206
rect 37740 585142 37792 585148
rect 37752 516089 37780 585142
rect 37844 563718 37872 636239
rect 38474 635352 38530 635361
rect 38474 635287 38530 635296
rect 38014 632224 38070 632233
rect 38014 632159 38070 632168
rect 37924 596284 37976 596290
rect 37924 596226 37976 596232
rect 37832 563712 37884 563718
rect 37832 563654 37884 563660
rect 37844 517449 37872 563654
rect 37830 517440 37886 517449
rect 37830 517375 37886 517384
rect 37738 516080 37794 516089
rect 37738 516015 37794 516024
rect 37830 507920 37886 507929
rect 37830 507855 37886 507864
rect 37738 488336 37794 488345
rect 37738 488271 37794 488280
rect 37648 477352 37700 477358
rect 37648 477294 37700 477300
rect 37752 368393 37780 488271
rect 37844 479806 37872 507855
rect 37832 479800 37884 479806
rect 37832 479742 37884 479748
rect 37936 478446 37964 596226
rect 38028 513369 38056 632159
rect 38106 630728 38162 630737
rect 38106 630663 38162 630672
rect 38014 513360 38070 513369
rect 38014 513295 38070 513304
rect 38028 479874 38056 513295
rect 38120 511057 38148 630663
rect 38290 629368 38346 629377
rect 38290 629303 38346 629312
rect 38198 628008 38254 628017
rect 38198 627943 38254 627952
rect 38106 511048 38162 511057
rect 38106 510983 38162 510992
rect 38120 480078 38148 510983
rect 38212 507929 38240 627943
rect 38304 509969 38332 629303
rect 38384 596760 38436 596766
rect 38384 596702 38436 596708
rect 38290 509960 38346 509969
rect 38290 509895 38346 509904
rect 38198 507920 38254 507929
rect 38198 507855 38254 507864
rect 38108 480072 38160 480078
rect 38108 480014 38160 480020
rect 38304 480010 38332 509895
rect 38292 480004 38344 480010
rect 38292 479946 38344 479952
rect 38016 479868 38068 479874
rect 38016 479810 38068 479816
rect 37924 478440 37976 478446
rect 37924 478382 37976 478388
rect 38396 477154 38424 596702
rect 38488 585818 38516 635287
rect 38566 610056 38622 610065
rect 38566 609991 38622 610000
rect 38476 585812 38528 585818
rect 38476 585754 38528 585760
rect 38488 585206 38516 585754
rect 38476 585200 38528 585206
rect 38476 585142 38528 585148
rect 38474 514040 38530 514049
rect 38474 513975 38530 513984
rect 38488 480049 38516 513975
rect 38580 489977 38608 609991
rect 39960 599978 39988 683318
rect 39960 599950 40080 599978
rect 39854 597408 39910 597417
rect 39854 597343 39910 597352
rect 39212 597236 39264 597242
rect 39212 597178 39264 597184
rect 39120 596216 39172 596222
rect 39120 596158 39172 596164
rect 39028 563304 39080 563310
rect 39028 563246 39080 563252
rect 39040 499574 39068 563246
rect 38948 499546 39068 499574
rect 38566 489968 38622 489977
rect 38566 489903 38622 489912
rect 38474 480040 38530 480049
rect 38474 479975 38530 479984
rect 38580 479942 38608 489903
rect 38948 484974 38976 499546
rect 39028 485308 39080 485314
rect 39028 485250 39080 485256
rect 38936 484968 38988 484974
rect 38936 484910 38988 484916
rect 38568 479936 38620 479942
rect 38568 479878 38620 479884
rect 38384 477148 38436 477154
rect 38384 477090 38436 477096
rect 39040 476882 39068 485250
rect 39132 478922 39160 596158
rect 39120 478916 39172 478922
rect 39120 478858 39172 478864
rect 39224 478582 39252 597178
rect 39578 597136 39634 597145
rect 39578 597071 39634 597080
rect 39488 596896 39540 596902
rect 39488 596838 39540 596844
rect 39396 596692 39448 596698
rect 39396 596634 39448 596640
rect 39304 596624 39356 596630
rect 39304 596566 39356 596572
rect 39212 478576 39264 478582
rect 39212 478518 39264 478524
rect 39316 477290 39344 596566
rect 39304 477284 39356 477290
rect 39304 477226 39356 477232
rect 39408 477222 39436 596634
rect 39396 477216 39448 477222
rect 39396 477158 39448 477164
rect 39500 477018 39528 596838
rect 39488 477012 39540 477018
rect 39488 476954 39540 476960
rect 39592 476950 39620 597071
rect 39672 596964 39724 596970
rect 39672 596906 39724 596912
rect 39684 485314 39712 596906
rect 39764 596828 39816 596834
rect 39764 596770 39816 596776
rect 39776 485314 39804 596770
rect 39672 485308 39724 485314
rect 39672 485250 39724 485256
rect 39764 485308 39816 485314
rect 39764 485250 39816 485256
rect 39868 485194 39896 597343
rect 39948 597032 40000 597038
rect 39948 596974 40000 596980
rect 39684 485166 39896 485194
rect 39580 476944 39632 476950
rect 39580 476886 39632 476892
rect 39028 476876 39080 476882
rect 39028 476818 39080 476824
rect 39684 476814 39712 485166
rect 39764 485104 39816 485110
rect 39960 485058 39988 596974
rect 40052 563310 40080 599950
rect 56414 597544 56470 597553
rect 56414 597479 56470 597488
rect 63222 597544 63278 597553
rect 63222 597479 63278 597488
rect 64234 597544 64290 597553
rect 64234 597479 64290 597488
rect 64878 597544 64934 597553
rect 64878 597479 64934 597488
rect 66810 597544 66866 597553
rect 66810 597479 66812 597488
rect 56428 597145 56456 597479
rect 56414 597136 56470 597145
rect 56414 597071 56470 597080
rect 56598 597136 56654 597145
rect 56598 597071 56654 597080
rect 59358 597136 59414 597145
rect 59358 597071 59414 597080
rect 56612 597038 56640 597071
rect 56600 597032 56652 597038
rect 56600 596974 56652 596980
rect 59372 596970 59400 597071
rect 59360 596964 59412 596970
rect 59360 596906 59412 596912
rect 63236 596902 63264 597479
rect 63224 596896 63276 596902
rect 63224 596838 63276 596844
rect 64248 596834 64276 597479
rect 64236 596828 64288 596834
rect 64236 596770 64288 596776
rect 64892 596766 64920 597479
rect 66864 597479 66866 597488
rect 67638 597544 67694 597553
rect 67638 597479 67694 597488
rect 68926 597544 68982 597553
rect 68926 597479 68982 597488
rect 69754 597544 69810 597553
rect 69754 597479 69810 597488
rect 71686 597544 71742 597553
rect 71686 597479 71742 597488
rect 73158 597544 73214 597553
rect 73158 597479 73214 597488
rect 74446 597544 74502 597553
rect 74446 597479 74502 597488
rect 74906 597544 74962 597553
rect 74906 597479 74962 597488
rect 77206 597544 77262 597553
rect 77206 597479 77262 597488
rect 78034 597544 78090 597553
rect 78034 597479 78090 597488
rect 78586 597544 78642 597553
rect 78586 597479 78642 597488
rect 81346 597544 81402 597553
rect 81346 597479 81402 597488
rect 84198 597544 84254 597553
rect 84198 597479 84200 597488
rect 66812 597450 66864 597456
rect 66168 597304 66220 597310
rect 66168 597246 66220 597252
rect 66180 596766 66208 597246
rect 64880 596760 64932 596766
rect 55402 596728 55458 596737
rect 64880 596702 64932 596708
rect 66168 596760 66220 596766
rect 66168 596702 66220 596708
rect 66824 596698 66852 597450
rect 55402 596663 55458 596672
rect 66812 596692 66864 596698
rect 55416 596222 55444 596663
rect 66812 596634 66864 596640
rect 67652 596562 67680 597479
rect 68834 597408 68890 597417
rect 68744 597372 68796 597378
rect 68834 597343 68890 597352
rect 68744 597314 68796 597320
rect 68756 596562 68784 597314
rect 68848 597174 68876 597343
rect 68836 597168 68888 597174
rect 68836 597110 68888 597116
rect 68848 596630 68876 597110
rect 68836 596624 68888 596630
rect 68836 596566 68888 596572
rect 67640 596556 67692 596562
rect 67640 596498 67692 596504
rect 68744 596556 68796 596562
rect 68744 596498 68796 596504
rect 55404 596216 55456 596222
rect 55404 596158 55456 596164
rect 68940 565049 68968 597479
rect 69768 597038 69796 597479
rect 71318 597408 71374 597417
rect 71318 597343 71374 597352
rect 69756 597032 69808 597038
rect 69756 596974 69808 596980
rect 69768 596494 69796 596974
rect 71332 596970 71360 597343
rect 70400 596964 70452 596970
rect 70400 596906 70452 596912
rect 71320 596964 71372 596970
rect 71320 596906 71372 596912
rect 69756 596488 69808 596494
rect 69756 596430 69808 596436
rect 70412 596426 70440 596906
rect 70400 596420 70452 596426
rect 70400 596362 70452 596368
rect 71700 566409 71728 597479
rect 71778 597408 71834 597417
rect 71778 597343 71834 597352
rect 71792 596426 71820 597343
rect 71780 596420 71832 596426
rect 71780 596362 71832 596368
rect 71792 594250 71820 596362
rect 73172 596358 73200 597479
rect 73160 596352 73212 596358
rect 73160 596294 73212 596300
rect 71780 594244 71832 594250
rect 71780 594186 71832 594192
rect 73172 594182 73200 596294
rect 73160 594176 73212 594182
rect 73160 594118 73212 594124
rect 74460 570761 74488 597479
rect 74920 597446 74948 597479
rect 74908 597440 74960 597446
rect 74908 597382 74960 597388
rect 76010 597408 76066 597417
rect 74920 597242 74948 597382
rect 76010 597343 76066 597352
rect 77114 597408 77170 597417
rect 77114 597343 77170 597352
rect 74908 597236 74960 597242
rect 74908 597178 74960 597184
rect 76024 596494 76052 597343
rect 77128 597242 77156 597343
rect 77116 597236 77168 597242
rect 77116 597178 77168 597184
rect 76012 596488 76064 596494
rect 76012 596430 76064 596436
rect 76024 594114 76052 596430
rect 77128 596290 77156 597178
rect 77116 596284 77168 596290
rect 77116 596226 77168 596232
rect 76012 594108 76064 594114
rect 76012 594050 76064 594056
rect 74446 570752 74502 570761
rect 74446 570687 74502 570696
rect 71686 566400 71742 566409
rect 71686 566335 71742 566344
rect 77220 565146 77248 597479
rect 78048 597106 78076 597479
rect 78036 597100 78088 597106
rect 78036 597042 78088 597048
rect 78600 565214 78628 597479
rect 81360 565282 81388 597479
rect 84252 597479 84254 597488
rect 86866 597544 86922 597553
rect 86866 597479 86922 597488
rect 88246 597544 88302 597553
rect 88246 597479 88302 597488
rect 92478 597544 92534 597553
rect 92478 597479 92534 597488
rect 93766 597544 93822 597553
rect 93766 597479 93822 597488
rect 124126 597544 124182 597553
rect 124126 597479 124182 597488
rect 129646 597544 129702 597553
rect 129646 597479 129702 597488
rect 131026 597544 131082 597553
rect 131026 597479 131082 597488
rect 133786 597544 133842 597553
rect 133786 597479 133842 597488
rect 136546 597544 136602 597553
rect 136546 597479 136602 597488
rect 142066 597544 142122 597553
rect 142066 597479 142122 597488
rect 146206 597544 146262 597553
rect 146206 597479 146262 597488
rect 84200 597450 84252 597456
rect 82818 597408 82874 597417
rect 82818 597343 82874 597352
rect 85580 597372 85632 597378
rect 82832 597310 82860 597343
rect 85580 597314 85632 597320
rect 82820 597304 82872 597310
rect 81438 597272 81494 597281
rect 85592 597281 85620 597314
rect 82820 597246 82872 597252
rect 85578 597272 85634 597281
rect 81438 597207 81494 597216
rect 85578 597207 85634 597216
rect 81452 596902 81480 597207
rect 81440 596896 81492 596902
rect 81440 596838 81492 596844
rect 82818 596864 82874 596873
rect 82818 596799 82820 596808
rect 82872 596799 82874 596808
rect 82820 596770 82872 596776
rect 84106 596456 84162 596465
rect 84106 596391 84162 596400
rect 84120 565350 84148 596391
rect 86880 565418 86908 597479
rect 86958 597272 87014 597281
rect 86958 597207 87014 597216
rect 86972 597174 87000 597207
rect 86960 597168 87012 597174
rect 86960 597110 87012 597116
rect 88260 565486 88288 597479
rect 92492 597446 92520 597479
rect 92480 597440 92532 597446
rect 92480 597382 92532 597388
rect 88338 597136 88394 597145
rect 88338 597071 88394 597080
rect 89718 597136 89774 597145
rect 89718 597071 89774 597080
rect 88352 597038 88380 597071
rect 88340 597032 88392 597038
rect 88340 596974 88392 596980
rect 89732 596970 89760 597071
rect 89720 596964 89772 596970
rect 89720 596906 89772 596912
rect 91190 596592 91246 596601
rect 91190 596527 91246 596536
rect 91098 596456 91154 596465
rect 91098 596391 91100 596400
rect 91152 596391 91154 596400
rect 91100 596362 91152 596368
rect 91204 596358 91232 596527
rect 91192 596352 91244 596358
rect 91006 596320 91062 596329
rect 91192 596294 91244 596300
rect 91006 596255 91062 596264
rect 91020 596222 91048 596255
rect 91008 596216 91060 596222
rect 91008 596158 91060 596164
rect 88248 565480 88300 565486
rect 88248 565422 88300 565428
rect 86868 565412 86920 565418
rect 86868 565354 86920 565360
rect 84108 565344 84160 565350
rect 84108 565286 84160 565292
rect 81348 565276 81400 565282
rect 81348 565218 81400 565224
rect 78588 565208 78640 565214
rect 93780 565185 93808 597479
rect 108946 597408 109002 597417
rect 108946 597343 109002 597352
rect 117226 597408 117282 597417
rect 117226 597343 117282 597352
rect 121366 597408 121422 597417
rect 121366 597343 121422 597352
rect 95238 597272 95294 597281
rect 95238 597207 95240 597216
rect 95292 597207 95294 597216
rect 95240 597178 95292 597184
rect 96618 597136 96674 597145
rect 96618 597071 96620 597080
rect 96672 597071 96674 597080
rect 96620 597042 96672 597048
rect 102046 596728 102102 596737
rect 102046 596663 102102 596672
rect 94042 596592 94098 596601
rect 94042 596527 94098 596536
rect 94056 596494 94084 596527
rect 94044 596488 94096 596494
rect 94044 596430 94096 596436
rect 96526 596456 96582 596465
rect 96526 596391 96582 596400
rect 99286 596456 99342 596465
rect 102060 596426 102088 596663
rect 106186 596592 106242 596601
rect 108960 596562 108988 597343
rect 114466 597272 114522 597281
rect 114466 597207 114522 597216
rect 111706 597000 111762 597009
rect 111706 596935 111762 596944
rect 111720 596698 111748 596935
rect 114480 596766 114508 597207
rect 117240 596834 117268 597343
rect 118606 597000 118662 597009
rect 118606 596935 118608 596944
rect 118660 596935 118662 596944
rect 118608 596906 118660 596912
rect 121380 596902 121408 597343
rect 121368 596896 121420 596902
rect 121368 596838 121420 596844
rect 117228 596828 117280 596834
rect 117228 596770 117280 596776
rect 114468 596760 114520 596766
rect 114468 596702 114520 596708
rect 111708 596692 111760 596698
rect 111708 596634 111760 596640
rect 124140 596630 124168 597479
rect 126886 597136 126942 597145
rect 126886 597071 126942 597080
rect 126900 597038 126928 597071
rect 126888 597032 126940 597038
rect 126888 596974 126940 596980
rect 124128 596624 124180 596630
rect 124128 596566 124180 596572
rect 106186 596527 106242 596536
rect 108948 596556 109000 596562
rect 106200 596494 106228 596527
rect 108948 596498 109000 596504
rect 106188 596488 106240 596494
rect 106188 596430 106240 596436
rect 99286 596391 99342 596400
rect 102048 596420 102100 596426
rect 96540 596290 96568 596391
rect 99300 596358 99328 596391
rect 102048 596362 102100 596368
rect 99288 596352 99340 596358
rect 99288 596294 99340 596300
rect 96528 596284 96580 596290
rect 96528 596226 96580 596232
rect 129660 565321 129688 597479
rect 131040 565554 131068 597479
rect 133800 565622 133828 597479
rect 136560 565690 136588 597479
rect 139306 597136 139362 597145
rect 139306 597071 139308 597080
rect 139360 597071 139362 597080
rect 139308 597042 139360 597048
rect 142080 565758 142108 597479
rect 142068 565752 142120 565758
rect 142068 565694 142120 565700
rect 136548 565684 136600 565690
rect 136548 565626 136600 565632
rect 133788 565616 133840 565622
rect 133788 565558 133840 565564
rect 131028 565548 131080 565554
rect 131028 565490 131080 565496
rect 146220 565457 146248 597479
rect 170864 567180 170916 567186
rect 170864 567122 170916 567128
rect 170876 565865 170904 567122
rect 170862 565856 170918 565865
rect 170862 565791 170918 565800
rect 146206 565448 146262 565457
rect 146206 565383 146262 565392
rect 129646 565312 129702 565321
rect 129646 565247 129702 565256
rect 78588 565150 78640 565156
rect 93766 565176 93822 565185
rect 77208 565140 77260 565146
rect 93766 565111 93822 565120
rect 77208 565082 77260 565088
rect 68926 565040 68982 565049
rect 68926 564975 68982 564984
rect 40040 563304 40092 563310
rect 40040 563246 40092 563252
rect 39764 485046 39816 485052
rect 39776 477086 39804 485046
rect 39868 485030 39988 485058
rect 39764 477080 39816 477086
rect 39764 477022 39816 477028
rect 39672 476808 39724 476814
rect 39672 476750 39724 476756
rect 39868 476746 39896 485030
rect 39948 484968 40000 484974
rect 39948 484910 40000 484916
rect 39960 480026 39988 484910
rect 39960 479998 40080 480026
rect 39856 476740 39908 476746
rect 39856 476682 39908 476688
rect 40052 443306 40080 479998
rect 56046 479632 56102 479641
rect 56046 479567 56102 479576
rect 56060 478922 56088 479567
rect 56048 478916 56100 478922
rect 56048 478858 56100 478864
rect 72330 478680 72386 478689
rect 74630 478680 74686 478689
rect 72330 478615 72332 478624
rect 72384 478615 72386 478624
rect 73804 478644 73856 478650
rect 72332 478586 72384 478592
rect 74630 478615 74686 478624
rect 73804 478586 73856 478592
rect 73158 478544 73214 478553
rect 73158 478479 73160 478488
rect 73212 478479 73214 478488
rect 73160 478450 73212 478456
rect 70860 477488 70912 477494
rect 63222 477456 63278 477465
rect 63222 477391 63278 477400
rect 64234 477456 64290 477465
rect 64234 477391 64290 477400
rect 64878 477456 64934 477465
rect 64878 477391 64934 477400
rect 66534 477456 66590 477465
rect 66534 477391 66590 477400
rect 67638 477456 67694 477465
rect 67638 477391 67694 477400
rect 68742 477456 68798 477465
rect 68742 477391 68798 477400
rect 70214 477456 70270 477465
rect 70214 477391 70216 477400
rect 59450 477320 59506 477329
rect 59450 477255 59506 477264
rect 60738 477320 60794 477329
rect 60738 477255 60794 477264
rect 58162 476912 58218 476921
rect 59464 476882 59492 477255
rect 60752 476950 60780 477255
rect 63236 477018 63264 477391
rect 63500 477080 63552 477086
rect 63500 477022 63552 477028
rect 63224 477012 63276 477018
rect 63224 476954 63276 476960
rect 60740 476944 60792 476950
rect 60740 476886 60792 476892
rect 58162 476847 58218 476856
rect 59452 476876 59504 476882
rect 58176 476814 58204 476847
rect 59452 476818 59504 476824
rect 63512 476814 63540 477022
rect 64248 476814 64276 477391
rect 64892 477154 64920 477391
rect 66548 477222 66576 477391
rect 67652 477358 67680 477391
rect 67640 477352 67692 477358
rect 67640 477294 67692 477300
rect 68756 477290 68784 477391
rect 70268 477391 70270 477400
rect 70858 477456 70860 477465
rect 70912 477456 70914 477465
rect 70858 477391 70914 477400
rect 70216 477362 70268 477368
rect 68744 477284 68796 477290
rect 68744 477226 68796 477232
rect 66536 477216 66588 477222
rect 66536 477158 66588 477164
rect 67548 477216 67600 477222
rect 67548 477158 67600 477164
rect 64880 477148 64932 477154
rect 64880 477090 64932 477096
rect 58164 476808 58216 476814
rect 57886 476776 57942 476785
rect 58164 476750 58216 476756
rect 63500 476808 63552 476814
rect 63500 476750 63552 476756
rect 64236 476808 64288 476814
rect 64236 476750 64288 476756
rect 64892 476746 64920 477090
rect 57886 476711 57888 476720
rect 57940 476711 57942 476720
rect 64880 476740 64932 476746
rect 57888 476682 57940 476688
rect 64880 476682 64932 476688
rect 67560 476678 67588 477158
rect 70228 476950 70256 477362
rect 70872 477018 70900 477391
rect 70860 477012 70912 477018
rect 70860 476954 70912 476960
rect 70216 476944 70268 476950
rect 70216 476886 70268 476892
rect 67548 476672 67600 476678
rect 67548 476614 67600 476620
rect 73172 476542 73200 478450
rect 73160 476536 73212 476542
rect 73160 476478 73212 476484
rect 73816 476474 73844 478586
rect 74644 478582 74672 478615
rect 74632 478576 74684 478582
rect 77208 478576 77260 478582
rect 74632 478518 74684 478524
rect 76930 478544 76986 478553
rect 77208 478518 77260 478524
rect 76930 478479 76986 478488
rect 76944 478446 76972 478479
rect 76932 478440 76984 478446
rect 75826 478408 75882 478417
rect 76932 478382 76984 478388
rect 75826 478343 75828 478352
rect 75880 478343 75882 478352
rect 75828 478314 75880 478320
rect 77220 477154 77248 478518
rect 78588 478440 78640 478446
rect 78588 478382 78640 478388
rect 78220 478372 78272 478378
rect 78220 478314 78272 478320
rect 78128 478304 78180 478310
rect 78128 478246 78180 478252
rect 78140 477465 78168 478246
rect 78126 477456 78182 477465
rect 78126 477391 78182 477400
rect 78140 477290 78168 477391
rect 78128 477284 78180 477290
rect 78128 477226 78180 477232
rect 77208 477148 77260 477154
rect 77208 477090 77260 477096
rect 78232 476610 78260 478314
rect 78600 477358 78628 478382
rect 79506 478272 79562 478281
rect 79506 478207 79508 478216
rect 79560 478207 79562 478216
rect 79508 478178 79560 478184
rect 80612 478168 80664 478174
rect 80610 478136 80612 478145
rect 82728 478168 82780 478174
rect 80664 478136 80666 478145
rect 82728 478110 82780 478116
rect 80610 478071 80666 478080
rect 81346 477456 81402 477465
rect 81346 477391 81402 477400
rect 81806 477456 81862 477465
rect 81806 477391 81862 477400
rect 78588 477352 78640 477358
rect 78588 477294 78640 477300
rect 78220 476604 78272 476610
rect 78220 476546 78272 476552
rect 73804 476468 73856 476474
rect 73804 476410 73856 476416
rect 68926 476232 68982 476241
rect 68926 476167 68982 476176
rect 71686 476232 71742 476241
rect 71686 476167 71742 476176
rect 74446 476232 74502 476241
rect 74446 476167 74502 476176
rect 77206 476232 77262 476241
rect 77206 476167 77262 476176
rect 78586 476232 78642 476241
rect 78586 476167 78642 476176
rect 68940 445058 68968 476167
rect 71700 449206 71728 476167
rect 71688 449200 71740 449206
rect 71688 449142 71740 449148
rect 68928 445052 68980 445058
rect 68928 444994 68980 445000
rect 74460 443601 74488 476167
rect 77220 443698 77248 476167
rect 78600 447846 78628 476167
rect 81360 447914 81388 477391
rect 81820 476882 81848 477391
rect 81808 476876 81860 476882
rect 81808 476818 81860 476824
rect 82636 476876 82688 476882
rect 82636 476818 82688 476824
rect 82648 476202 82676 476818
rect 82740 476241 82768 478110
rect 86314 477592 86370 477601
rect 86314 477527 86370 477536
rect 82818 477456 82874 477465
rect 82818 477391 82874 477400
rect 84106 477456 84162 477465
rect 84106 477391 84162 477400
rect 85302 477456 85358 477465
rect 86328 477426 86356 477527
rect 86960 477488 87012 477494
rect 86866 477456 86922 477465
rect 85302 477391 85358 477400
rect 85580 477420 85632 477426
rect 82832 476814 82860 477391
rect 82820 476808 82872 476814
rect 82820 476750 82872 476756
rect 83924 476808 83976 476814
rect 83924 476750 83976 476756
rect 82726 476232 82782 476241
rect 82636 476196 82688 476202
rect 82726 476167 82782 476176
rect 82636 476138 82688 476144
rect 83936 476134 83964 476750
rect 84016 476740 84068 476746
rect 84016 476682 84068 476688
rect 84028 476649 84056 476682
rect 84014 476640 84070 476649
rect 84014 476575 84070 476584
rect 84028 476338 84056 476575
rect 84016 476332 84068 476338
rect 84016 476274 84068 476280
rect 83924 476128 83976 476134
rect 83924 476070 83976 476076
rect 84120 447982 84148 477391
rect 85316 476678 85344 477391
rect 85580 477362 85632 477368
rect 86316 477420 86368 477426
rect 87604 477488 87656 477494
rect 86960 477430 87012 477436
rect 87602 477456 87604 477465
rect 87656 477456 87658 477465
rect 86866 477391 86922 477400
rect 86316 477362 86368 477368
rect 85592 477222 85620 477362
rect 85580 477216 85632 477222
rect 85580 477158 85632 477164
rect 85304 476672 85356 476678
rect 85304 476614 85356 476620
rect 86880 448050 86908 477391
rect 86972 477086 87000 477430
rect 87602 477391 87658 477400
rect 88246 477456 88302 477465
rect 88246 477391 88302 477400
rect 88706 477456 88762 477465
rect 88706 477391 88762 477400
rect 89718 477456 89774 477465
rect 89718 477391 89774 477400
rect 91190 477456 91246 477465
rect 91190 477391 91246 477400
rect 92202 477456 92258 477465
rect 92202 477391 92258 477400
rect 93030 477456 93086 477465
rect 93030 477391 93086 477400
rect 94410 477456 94466 477465
rect 94410 477391 94466 477400
rect 95790 477456 95846 477465
rect 95790 477391 95846 477400
rect 96986 477456 97042 477465
rect 96986 477391 97042 477400
rect 86960 477080 87012 477086
rect 86960 477022 87012 477028
rect 88260 448118 88288 477391
rect 88720 476950 88748 477391
rect 89732 477018 89760 477391
rect 89720 477012 89772 477018
rect 89720 476954 89772 476960
rect 88708 476944 88760 476950
rect 88708 476886 88760 476892
rect 89732 476814 89760 476954
rect 91100 476944 91152 476950
rect 91100 476886 91152 476892
rect 89720 476808 89772 476814
rect 89720 476750 89772 476756
rect 91112 476542 91140 476886
rect 91100 476536 91152 476542
rect 91006 476504 91062 476513
rect 91100 476478 91152 476484
rect 91006 476439 91062 476448
rect 91020 448186 91048 476439
rect 91204 476406 91232 477391
rect 92216 476950 92244 477391
rect 93044 477154 93072 477391
rect 93032 477148 93084 477154
rect 93032 477090 93084 477096
rect 92204 476944 92256 476950
rect 92204 476886 92256 476892
rect 91284 476672 91336 476678
rect 91284 476614 91336 476620
rect 91192 476400 91244 476406
rect 91192 476342 91244 476348
rect 91204 476270 91232 476342
rect 91296 476270 91324 476614
rect 93044 476542 93072 477090
rect 93032 476536 93084 476542
rect 93032 476478 93084 476484
rect 93766 476504 93822 476513
rect 94424 476474 94452 477391
rect 95804 477358 95832 477391
rect 95792 477352 95844 477358
rect 95792 477294 95844 477300
rect 96528 477352 96580 477358
rect 96528 477294 96580 477300
rect 96540 477086 96568 477294
rect 97000 477290 97028 477391
rect 96988 477284 97040 477290
rect 96988 477226 97040 477232
rect 96528 477080 96580 477086
rect 96528 477022 96580 477028
rect 95974 476504 96030 476513
rect 93766 476439 93822 476448
rect 94412 476468 94464 476474
rect 91192 476264 91244 476270
rect 91192 476206 91244 476212
rect 91284 476264 91336 476270
rect 91284 476206 91336 476212
rect 91008 448180 91060 448186
rect 91008 448122 91060 448128
rect 88248 448112 88300 448118
rect 88248 448054 88300 448060
rect 86868 448044 86920 448050
rect 86868 447986 86920 447992
rect 84108 447976 84160 447982
rect 84108 447918 84160 447924
rect 81348 447908 81400 447914
rect 81348 447850 81400 447856
rect 78588 447840 78640 447846
rect 78588 447782 78640 447788
rect 93780 444961 93808 476439
rect 95974 476439 96030 476448
rect 94412 476410 94464 476416
rect 95988 476241 96016 476439
rect 95974 476232 96030 476241
rect 95974 476167 96030 476176
rect 96526 476232 96582 476241
rect 96526 476167 96582 476176
rect 99286 476232 99342 476241
rect 99286 476167 99342 476176
rect 102046 476232 102102 476241
rect 102046 476167 102102 476176
rect 104806 476232 104862 476241
rect 104806 476167 104862 476176
rect 106186 476232 106242 476241
rect 106186 476167 106242 476176
rect 108946 476232 109002 476241
rect 108946 476167 109002 476176
rect 111706 476232 111762 476241
rect 111706 476167 111762 476176
rect 114466 476232 114522 476241
rect 114466 476167 114522 476176
rect 117226 476232 117282 476241
rect 117226 476167 117282 476176
rect 118606 476232 118662 476241
rect 118606 476167 118662 476176
rect 121366 476232 121422 476241
rect 121366 476167 121422 476176
rect 124126 476232 124182 476241
rect 124126 476167 124182 476176
rect 126886 476232 126942 476241
rect 126886 476167 126942 476176
rect 129646 476232 129702 476241
rect 129646 476167 129702 476176
rect 131026 476232 131082 476241
rect 131026 476167 131082 476176
rect 133786 476232 133842 476241
rect 133786 476167 133842 476176
rect 136546 476232 136602 476241
rect 136546 476167 136602 476176
rect 139306 476232 139362 476241
rect 139306 476167 139362 476176
rect 142066 476232 142122 476241
rect 142066 476167 142122 476176
rect 143446 476232 143502 476241
rect 143446 476167 143502 476176
rect 146206 476232 146262 476241
rect 146206 476167 146262 476176
rect 96540 445126 96568 476167
rect 99300 445194 99328 476167
rect 102060 445262 102088 476167
rect 104820 445330 104848 476167
rect 106200 445398 106228 476167
rect 106188 445392 106240 445398
rect 106188 445334 106240 445340
rect 104808 445324 104860 445330
rect 104808 445266 104860 445272
rect 102048 445256 102100 445262
rect 102048 445198 102100 445204
rect 99288 445188 99340 445194
rect 99288 445130 99340 445136
rect 96528 445120 96580 445126
rect 108960 445097 108988 476167
rect 111720 445233 111748 476167
rect 114480 445466 114508 476167
rect 117240 445534 117268 476167
rect 118620 445602 118648 476167
rect 121380 445670 121408 476167
rect 124140 445738 124168 476167
rect 124128 445732 124180 445738
rect 124128 445674 124180 445680
rect 121368 445664 121420 445670
rect 121368 445606 121420 445612
rect 118608 445596 118660 445602
rect 118608 445538 118660 445544
rect 117228 445528 117280 445534
rect 117228 445470 117280 445476
rect 114468 445460 114520 445466
rect 114468 445402 114520 445408
rect 111706 445224 111762 445233
rect 111706 445159 111762 445168
rect 96528 445062 96580 445068
rect 108946 445088 109002 445097
rect 108946 445023 109002 445032
rect 126900 444990 126928 476167
rect 126888 444984 126940 444990
rect 93766 444952 93822 444961
rect 126888 444926 126940 444932
rect 129660 444922 129688 476167
rect 131040 448254 131068 476167
rect 133800 448322 133828 476167
rect 136560 448390 136588 476167
rect 139320 448458 139348 476167
rect 142080 448526 142108 476167
rect 142068 448520 142120 448526
rect 142068 448462 142120 448468
rect 139308 448452 139360 448458
rect 139308 448394 139360 448400
rect 136548 448384 136600 448390
rect 136548 448326 136600 448332
rect 133788 448316 133840 448322
rect 133788 448258 133840 448264
rect 131028 448248 131080 448254
rect 131028 448190 131080 448196
rect 143460 447778 143488 476167
rect 143448 447772 143500 447778
rect 143448 447714 143500 447720
rect 146220 447710 146248 476167
rect 146208 447704 146260 447710
rect 146208 447646 146260 447652
rect 170864 447092 170916 447098
rect 170864 447034 170916 447040
rect 170876 445777 170904 447034
rect 170862 445768 170918 445777
rect 170862 445703 170918 445712
rect 93766 444887 93822 444896
rect 129648 444916 129700 444922
rect 129648 444858 129700 444864
rect 77208 443692 77260 443698
rect 77208 443634 77260 443640
rect 74446 443592 74502 443601
rect 74446 443527 74502 443536
rect 38476 443284 38528 443290
rect 38476 443226 38528 443232
rect 39960 443278 40080 443306
rect 38488 397361 38516 443226
rect 38474 397352 38530 397361
rect 38474 397287 38530 397296
rect 38474 395448 38530 395457
rect 38474 395383 38530 395392
rect 37738 368384 37794 368393
rect 37738 368319 37794 368328
rect 38198 368384 38254 368393
rect 38198 368319 38254 368328
rect 38212 360058 38240 368319
rect 38382 367568 38438 367577
rect 38382 367503 38438 367512
rect 38200 360052 38252 360058
rect 38200 359994 38252 360000
rect 36544 357468 36596 357474
rect 36544 357410 36596 357416
rect 36556 340338 36584 357410
rect 38396 351218 38424 367503
rect 38488 358086 38516 395383
rect 39026 393544 39082 393553
rect 39026 393479 39082 393488
rect 38842 392320 38898 392329
rect 38842 392255 38898 392264
rect 38750 389464 38806 389473
rect 38750 389399 38806 389408
rect 38658 387832 38714 387841
rect 38658 387767 38714 387776
rect 38566 369880 38622 369889
rect 38566 369815 38622 369824
rect 38476 358080 38528 358086
rect 38476 358022 38528 358028
rect 38384 351212 38436 351218
rect 38384 351154 38436 351160
rect 38580 342922 38608 369815
rect 38568 342916 38620 342922
rect 38568 342858 38620 342864
rect 36544 340332 36596 340338
rect 36544 340274 36596 340280
rect 35164 308508 35216 308514
rect 35164 308450 35216 308456
rect 26884 301504 26936 301510
rect 26884 301446 26936 301452
rect 25504 298784 25556 298790
rect 25504 298726 25556 298732
rect 38672 296002 38700 387767
rect 38764 297430 38792 389399
rect 38856 354006 38884 392255
rect 38934 390688 38990 390697
rect 38934 390623 38990 390632
rect 38844 354000 38896 354006
rect 38844 353942 38896 353948
rect 38948 352578 38976 390623
rect 39040 355366 39068 393479
rect 39960 360074 39988 443278
rect 39960 360046 40080 360074
rect 39028 355360 39080 355366
rect 39028 355302 39080 355308
rect 38936 352572 38988 352578
rect 38936 352514 38988 352520
rect 38752 297424 38804 297430
rect 38752 297366 38804 297372
rect 38660 295996 38712 296002
rect 38660 295938 38712 295944
rect 40052 285054 40080 360046
rect 147588 358284 147640 358290
rect 147588 358226 147640 358232
rect 146852 358216 146904 358222
rect 61382 358184 61438 358193
rect 61382 358119 61438 358128
rect 64326 358184 64382 358193
rect 146852 358158 146904 358164
rect 64326 358119 64382 358128
rect 146484 358148 146536 358154
rect 56506 357368 56562 357377
rect 56506 357303 56562 357312
rect 59266 357368 59322 357377
rect 59266 357303 59322 357312
rect 60646 357368 60702 357377
rect 60646 357303 60702 357312
rect 56520 291854 56548 357303
rect 58622 357232 58678 357241
rect 58622 357167 58678 357176
rect 58636 294642 58664 357167
rect 59280 326466 59308 357303
rect 60660 356658 60688 357303
rect 60648 356652 60700 356658
rect 60648 356594 60700 356600
rect 61396 337414 61424 358119
rect 62026 357368 62082 357377
rect 62026 357303 62082 357312
rect 63406 357368 63462 357377
rect 63406 357303 63462 357312
rect 61384 337408 61436 337414
rect 61384 337350 61436 337356
rect 59268 326460 59320 326466
rect 59268 326402 59320 326408
rect 62040 316742 62068 357303
rect 62764 356652 62816 356658
rect 62764 356594 62816 356600
rect 62028 316736 62080 316742
rect 62028 316678 62080 316684
rect 62776 312594 62804 356594
rect 63420 330682 63448 357303
rect 64340 356114 64368 358119
rect 146484 358090 146536 358096
rect 67546 357368 67602 357377
rect 67546 357303 67602 357312
rect 68834 357368 68890 357377
rect 68834 357303 68890 357312
rect 70306 357368 70362 357377
rect 70306 357303 70362 357312
rect 71686 357368 71742 357377
rect 71686 357303 71742 357312
rect 73066 357368 73122 357377
rect 73066 357303 73122 357312
rect 74354 357368 74410 357377
rect 74354 357303 74410 357312
rect 75826 357368 75882 357377
rect 75826 357303 75882 357312
rect 76010 357368 76066 357377
rect 76010 357303 76066 357312
rect 78586 357368 78642 357377
rect 78586 357303 78642 357312
rect 79966 357368 80022 357377
rect 79966 357303 80022 357312
rect 81346 357368 81402 357377
rect 81346 357303 81402 357312
rect 86866 357368 86922 357377
rect 86866 357303 86922 357312
rect 88246 357368 88302 357377
rect 88246 357303 88302 357312
rect 91006 357368 91062 357377
rect 91006 357303 91062 357312
rect 93398 357368 93454 357377
rect 93398 357303 93454 357312
rect 96526 357368 96582 357377
rect 96526 357303 96582 357312
rect 99286 357368 99342 357377
rect 99286 357303 99342 357312
rect 102046 357368 102102 357377
rect 102046 357303 102102 357312
rect 106186 357368 106242 357377
rect 106186 357303 106242 357312
rect 66166 356144 66222 356153
rect 64328 356108 64380 356114
rect 64328 356050 64380 356056
rect 65524 356108 65576 356114
rect 66166 356079 66222 356088
rect 65524 356050 65576 356056
rect 63408 330676 63460 330682
rect 63408 330618 63460 330624
rect 65536 322318 65564 356050
rect 66180 323610 66208 356079
rect 66168 323604 66220 323610
rect 66168 323546 66220 323552
rect 65524 322312 65576 322318
rect 65524 322254 65576 322260
rect 62764 312588 62816 312594
rect 62764 312530 62816 312536
rect 67560 294710 67588 357303
rect 68848 327894 68876 357303
rect 68926 357096 68982 357105
rect 68926 357031 68982 357040
rect 68940 356250 68968 357031
rect 68928 356244 68980 356250
rect 68928 356186 68980 356192
rect 68926 356144 68982 356153
rect 68926 356079 68928 356088
rect 68980 356079 68982 356088
rect 68928 356050 68980 356056
rect 70320 329186 70348 357303
rect 71594 357232 71650 357241
rect 71594 357167 71650 357176
rect 70308 329180 70360 329186
rect 70308 329122 70360 329128
rect 68836 327888 68888 327894
rect 68836 327830 68888 327836
rect 71608 298858 71636 357167
rect 71596 298852 71648 298858
rect 71596 298794 71648 298800
rect 71700 296138 71728 357303
rect 73080 344418 73108 357303
rect 74078 357232 74134 357241
rect 74078 357167 74134 357176
rect 74092 356182 74120 357167
rect 74080 356176 74132 356182
rect 74080 356118 74132 356124
rect 73068 344412 73120 344418
rect 73068 344354 73120 344360
rect 74368 308446 74396 357303
rect 75840 318170 75868 357303
rect 76024 348566 76052 357303
rect 77022 357232 77078 357241
rect 77022 357167 77078 357176
rect 78494 357232 78550 357241
rect 78494 357167 78550 357176
rect 76012 348560 76064 348566
rect 76012 348502 76064 348508
rect 77036 340270 77064 357167
rect 77206 356416 77262 356425
rect 77206 356351 77262 356360
rect 77220 356318 77248 356351
rect 77208 356312 77260 356318
rect 77208 356254 77260 356260
rect 78508 347138 78536 357167
rect 78496 347132 78548 347138
rect 78496 347074 78548 347080
rect 77024 340264 77076 340270
rect 77024 340206 77076 340212
rect 75828 318164 75880 318170
rect 75828 318106 75880 318112
rect 78600 311234 78628 357303
rect 79980 320958 80008 357303
rect 81254 357232 81310 357241
rect 81254 357167 81310 357176
rect 81268 341698 81296 357167
rect 81256 341692 81308 341698
rect 81256 341634 81308 341640
rect 79968 320952 80020 320958
rect 79968 320894 80020 320900
rect 78588 311228 78640 311234
rect 78588 311170 78640 311176
rect 81360 309874 81388 357303
rect 84106 356688 84162 356697
rect 84106 356623 84162 356632
rect 81348 309868 81400 309874
rect 81348 309810 81400 309816
rect 74356 308440 74408 308446
rect 74356 308382 74408 308388
rect 71688 296132 71740 296138
rect 71688 296074 71740 296080
rect 67548 294704 67600 294710
rect 67548 294646 67600 294652
rect 58624 294636 58676 294642
rect 58624 294578 58676 294584
rect 84120 291922 84148 356623
rect 86880 293350 86908 357303
rect 87604 318844 87656 318850
rect 87604 318786 87656 318792
rect 86868 293344 86920 293350
rect 86868 293286 86920 293292
rect 84108 291916 84160 291922
rect 84108 291858 84160 291864
rect 56508 291848 56560 291854
rect 56508 291790 56560 291796
rect 87616 287774 87644 318786
rect 88260 314022 88288 357303
rect 91020 315382 91048 357303
rect 93412 349858 93440 357303
rect 93400 349852 93452 349858
rect 93400 349794 93452 349800
rect 91008 315376 91060 315382
rect 91008 315318 91060 315324
rect 88248 314016 88300 314022
rect 88248 313958 88300 313964
rect 90364 305040 90416 305046
rect 90364 304982 90416 304988
rect 89720 292596 89772 292602
rect 89720 292538 89772 292544
rect 89732 290494 89760 292538
rect 89720 290488 89772 290494
rect 89720 290430 89772 290436
rect 90376 289270 90404 304982
rect 96540 300150 96568 357303
rect 99300 301578 99328 357303
rect 102060 303006 102088 357303
rect 104806 356144 104862 356153
rect 104806 356079 104862 356088
rect 104820 304298 104848 356079
rect 106200 307154 106228 357303
rect 144642 355328 144698 355337
rect 144642 355263 144698 355272
rect 138754 353968 138810 353977
rect 138754 353903 138810 353912
rect 134340 348424 134392 348430
rect 134340 348366 134392 348372
rect 133604 347064 133656 347070
rect 133604 347006 133656 347012
rect 133236 327752 133288 327758
rect 133236 327694 133288 327700
rect 131764 324352 131816 324358
rect 131764 324294 131816 324300
rect 106188 307148 106240 307154
rect 106188 307090 106240 307096
rect 104808 304292 104860 304298
rect 104808 304234 104860 304240
rect 102048 303000 102100 303006
rect 102048 302942 102100 302948
rect 99288 301572 99340 301578
rect 99288 301514 99340 301520
rect 96528 300144 96580 300150
rect 96528 300086 96580 300092
rect 131396 298172 131448 298178
rect 131396 298114 131448 298120
rect 90364 289264 90416 289270
rect 90364 289206 90416 289212
rect 87604 287768 87656 287774
rect 87604 287710 87656 287716
rect 40040 285048 40092 285054
rect 40040 284990 40092 284996
rect 18604 284980 18656 284986
rect 18604 284922 18656 284928
rect 130568 283824 130620 283830
rect 130568 283766 130620 283772
rect 116676 283484 116728 283490
rect 116676 283426 116728 283432
rect 90364 282532 90416 282538
rect 90364 282474 90416 282480
rect 15844 282124 15896 282130
rect 15844 282066 15896 282072
rect 3516 280968 3568 280974
rect 3516 280910 3568 280916
rect 3424 279540 3476 279546
rect 3424 279482 3476 279488
rect 3332 267708 3384 267714
rect 3332 267650 3384 267656
rect 3344 267209 3372 267650
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 2964 255264 3016 255270
rect 2964 255206 3016 255212
rect 2976 254153 3004 255206
rect 2962 254144 3018 254153
rect 2962 254079 3018 254088
rect 3332 241460 3384 241466
rect 3332 241402 3384 241408
rect 3344 241097 3372 241402
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3056 215280 3108 215286
rect 3056 215222 3108 215228
rect 3068 214985 3096 215222
rect 3054 214976 3110 214985
rect 3054 214911 3110 214920
rect 3332 189032 3384 189038
rect 3332 188974 3384 188980
rect 3344 188873 3372 188974
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3056 164212 3108 164218
rect 3056 164154 3108 164160
rect 3068 162897 3096 164154
rect 3054 162888 3110 162897
rect 3054 162823 3110 162832
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3332 137964 3384 137970
rect 3332 137906 3384 137912
rect 3344 136785 3372 137906
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3332 97980 3384 97986
rect 3332 97922 3384 97928
rect 3344 97617 3372 97922
rect 3330 97608 3386 97617
rect 3330 97543 3386 97552
rect 1400 78056 1452 78062
rect 1400 77998 1452 78004
rect 20 77988 72 77994
rect 20 77930 72 77936
rect 32 16574 60 77930
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 77998
rect 3436 32473 3464 279482
rect 3528 58585 3556 280910
rect 3792 280900 3844 280906
rect 3792 280842 3844 280848
rect 3700 280832 3752 280838
rect 3700 280774 3752 280780
rect 3608 280220 3660 280226
rect 3608 280162 3660 280168
rect 3620 71641 3648 280162
rect 3712 84697 3740 280774
rect 3804 201929 3832 280842
rect 3790 201920 3846 201929
rect 3790 201855 3846 201864
rect 3698 84688 3754 84697
rect 3698 84623 3754 84632
rect 3606 71632 3662 71641
rect 3606 71567 3662 71576
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 15856 20670 15884 282066
rect 90376 97986 90404 282474
rect 115296 280492 115348 280498
rect 115296 280434 115348 280440
rect 115204 280288 115256 280294
rect 115204 280230 115256 280236
rect 115216 150414 115244 280230
rect 115308 255270 115336 280434
rect 116584 280356 116636 280362
rect 116584 280298 116636 280304
rect 115296 255264 115348 255270
rect 115296 255206 115348 255212
rect 115204 150408 115256 150414
rect 115204 150350 115256 150356
rect 116596 137970 116624 280298
rect 116688 164218 116716 283426
rect 119528 283416 119580 283422
rect 119528 283358 119580 283364
rect 119436 281852 119488 281858
rect 119436 281794 119488 281800
rect 119344 280424 119396 280430
rect 119344 280366 119396 280372
rect 116676 164212 116728 164218
rect 116676 164154 116728 164160
rect 116584 137964 116636 137970
rect 116584 137906 116636 137912
rect 90364 97980 90416 97986
rect 90364 97922 90416 97928
rect 119356 45558 119384 280366
rect 119448 189038 119476 281794
rect 119540 215286 119568 283358
rect 126152 283348 126204 283354
rect 126152 283290 126204 283296
rect 125416 283212 125468 283218
rect 125416 283154 125468 283160
rect 120908 281988 120960 281994
rect 120908 281930 120960 281936
rect 119620 281920 119672 281926
rect 119620 281862 119672 281868
rect 119632 241466 119660 281862
rect 120816 281784 120868 281790
rect 120816 281726 120868 281732
rect 120724 281716 120776 281722
rect 120724 281658 120776 281664
rect 119620 241460 119672 241466
rect 119620 241402 119672 241408
rect 119528 215280 119580 215286
rect 119528 215222 119580 215228
rect 119436 189032 119488 189038
rect 119436 188974 119488 188980
rect 119344 45552 119396 45558
rect 119344 45494 119396 45500
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 15844 20664 15896 20670
rect 15844 20606 15896 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 120736 6866 120764 281658
rect 120828 111790 120856 281726
rect 120920 267714 120948 281930
rect 121276 281648 121328 281654
rect 121276 281590 121328 281596
rect 124588 281648 124640 281654
rect 124588 281590 124640 281596
rect 120908 267708 120960 267714
rect 120908 267650 120960 267656
rect 120816 111784 120868 111790
rect 120816 111726 120868 111732
rect 121288 46918 121316 281590
rect 121368 280152 121420 280158
rect 121368 280094 121420 280100
rect 124220 280152 124272 280158
rect 124220 280094 124272 280100
rect 121276 46912 121328 46918
rect 121276 46854 121328 46860
rect 121380 20670 121408 280094
rect 124232 279970 124260 280094
rect 124600 279970 124628 281590
rect 125428 279970 125456 283154
rect 125506 281752 125562 281761
rect 125506 281687 125562 281696
rect 124232 279942 124476 279970
rect 124600 279942 124844 279970
rect 125212 279942 125456 279970
rect 125520 279970 125548 281687
rect 126164 279970 126192 283290
rect 127256 283280 127308 283286
rect 127256 283222 127308 283228
rect 126520 283008 126572 283014
rect 126520 282950 126572 282956
rect 126532 279970 126560 282950
rect 126886 281888 126942 281897
rect 126886 281823 126942 281832
rect 126900 279970 126928 281823
rect 127268 279970 127296 283222
rect 128268 283144 128320 283150
rect 128268 283086 128320 283092
rect 127624 282328 127676 282334
rect 127624 282270 127676 282276
rect 127636 279970 127664 282270
rect 127760 280256 127816 280265
rect 127760 280191 127816 280200
rect 125520 279942 125580 279970
rect 125948 279942 126192 279970
rect 126316 279942 126560 279970
rect 126684 279942 126928 279970
rect 127052 279942 127296 279970
rect 127420 279942 127664 279970
rect 127774 279956 127802 280191
rect 128280 279970 128308 283086
rect 129464 283076 129516 283082
rect 129464 283018 129516 283024
rect 129096 282192 129148 282198
rect 129096 282134 129148 282140
rect 128726 281616 128782 281625
rect 128726 281551 128782 281560
rect 128740 279970 128768 281551
rect 129108 279970 129136 282134
rect 129476 279970 129504 283018
rect 130200 282260 130252 282266
rect 130200 282202 130252 282208
rect 129556 280696 129608 280702
rect 129556 280638 129608 280644
rect 128156 279942 128308 279970
rect 128524 279942 128768 279970
rect 128892 279942 129136 279970
rect 129260 279942 129504 279970
rect 129568 279970 129596 280638
rect 130212 279970 130240 282202
rect 130580 279970 130608 283766
rect 130936 281036 130988 281042
rect 130936 280978 130988 280984
rect 130948 279970 130976 280978
rect 131028 280764 131080 280770
rect 131028 280706 131080 280712
rect 129568 279942 129628 279970
rect 129996 279942 130240 279970
rect 130364 279942 130608 279970
rect 130732 279942 130976 279970
rect 131040 279970 131068 280706
rect 131408 279970 131436 298114
rect 131776 279970 131804 324294
rect 132132 311908 132184 311914
rect 132132 311850 132184 311856
rect 132144 279970 132172 311850
rect 132868 289128 132920 289134
rect 132868 289070 132920 289076
rect 132592 287836 132644 287842
rect 132592 287778 132644 287784
rect 132604 280242 132632 287778
rect 132558 280214 132632 280242
rect 131040 279942 131100 279970
rect 131408 279942 131468 279970
rect 131776 279942 131836 279970
rect 132144 279942 132204 279970
rect 132558 279956 132586 280214
rect 132880 279970 132908 289070
rect 133248 279970 133276 327694
rect 133616 279970 133644 347006
rect 133970 290456 134026 290465
rect 133970 290391 134026 290400
rect 133788 282056 133840 282062
rect 133788 281998 133840 282004
rect 133800 280974 133828 281998
rect 133788 280968 133840 280974
rect 133788 280910 133840 280916
rect 133984 279970 134012 290391
rect 134352 279970 134380 348366
rect 136916 344344 136968 344350
rect 136916 344286 136968 344292
rect 135076 320884 135128 320890
rect 135076 320826 135128 320832
rect 134984 285184 135036 285190
rect 134984 285126 135036 285132
rect 134996 279970 135024 285126
rect 132880 279942 132940 279970
rect 133248 279942 133308 279970
rect 133616 279942 133676 279970
rect 133984 279942 134044 279970
rect 134352 279942 134412 279970
rect 134780 279942 135024 279970
rect 135088 279970 135116 320826
rect 136548 315308 136600 315314
rect 136548 315250 136600 315256
rect 135444 292120 135496 292126
rect 135444 292062 135496 292068
rect 135456 279970 135484 292062
rect 136454 284880 136510 284889
rect 136454 284815 136510 284824
rect 136088 283620 136140 283626
rect 136088 283562 136140 283568
rect 136100 279970 136128 283562
rect 136468 279970 136496 284815
rect 135088 279942 135148 279970
rect 135456 279942 135516 279970
rect 135884 279942 136128 279970
rect 136252 279942 136496 279970
rect 136560 279970 136588 315250
rect 136928 279970 136956 344286
rect 138020 326392 138072 326398
rect 138020 326334 138072 326340
rect 137652 323740 137704 323746
rect 137652 323682 137704 323688
rect 137284 305652 137336 305658
rect 137284 305594 137336 305600
rect 137296 279970 137324 305594
rect 137664 279970 137692 323682
rect 138032 279970 138060 326334
rect 138388 322244 138440 322250
rect 138388 322186 138440 322192
rect 138400 279970 138428 322186
rect 138768 279970 138796 353903
rect 142802 352608 142858 352617
rect 142802 352543 142858 352552
rect 141330 351112 141386 351121
rect 141330 351047 141386 351056
rect 140594 349752 140650 349761
rect 140594 349687 140650 349696
rect 140228 345704 140280 345710
rect 140228 345646 140280 345652
rect 139124 340196 139176 340202
rect 139124 340138 139176 340144
rect 139136 279970 139164 340138
rect 139860 338768 139912 338774
rect 139860 338710 139912 338716
rect 139492 318232 139544 318238
rect 139492 318174 139544 318180
rect 139504 279970 139532 318174
rect 139872 279970 139900 338710
rect 140240 279970 140268 345646
rect 140608 279970 140636 349687
rect 140962 290592 141018 290601
rect 140962 290527 141018 290536
rect 140976 279970 141004 290527
rect 141344 279970 141372 351047
rect 142436 341556 142488 341562
rect 142436 341498 142488 341504
rect 141700 333260 141752 333266
rect 141700 333202 141752 333208
rect 141712 279970 141740 333202
rect 142068 319456 142120 319462
rect 142068 319398 142120 319404
rect 142080 279970 142108 319398
rect 142448 279970 142476 341498
rect 142816 279970 142844 352543
rect 143906 337376 143962 337385
rect 143906 337311 143962 337320
rect 143540 330540 143592 330546
rect 143540 330482 143592 330488
rect 143172 324964 143224 324970
rect 143172 324906 143224 324912
rect 143184 279970 143212 324906
rect 143448 282940 143500 282946
rect 143448 282882 143500 282888
rect 143460 282334 143488 282882
rect 143448 282328 143500 282334
rect 143448 282270 143500 282276
rect 143448 281580 143500 281586
rect 143448 281522 143500 281528
rect 143460 280906 143488 281522
rect 143448 280900 143500 280906
rect 143448 280842 143500 280848
rect 143552 279970 143580 330482
rect 143920 279970 143948 337311
rect 144552 285252 144604 285258
rect 144552 285194 144604 285200
rect 144564 279970 144592 285194
rect 136560 279942 136620 279970
rect 136928 279942 136988 279970
rect 137296 279942 137356 279970
rect 137664 279942 137724 279970
rect 138032 279942 138092 279970
rect 138400 279942 138460 279970
rect 138768 279942 138828 279970
rect 139136 279942 139196 279970
rect 139504 279942 139564 279970
rect 139872 279942 139932 279970
rect 140240 279942 140300 279970
rect 140608 279942 140668 279970
rect 140976 279942 141036 279970
rect 141344 279942 141404 279970
rect 141712 279942 141772 279970
rect 142080 279942 142140 279970
rect 142448 279942 142508 279970
rect 142816 279942 142876 279970
rect 143184 279942 143244 279970
rect 143552 279942 143612 279970
rect 143920 279942 143980 279970
rect 144348 279942 144592 279970
rect 144656 279970 144684 355263
rect 145010 342952 145066 342961
rect 145010 342887 145066 342896
rect 145024 279970 145052 342887
rect 145746 327720 145802 327729
rect 145746 327655 145802 327664
rect 145656 285320 145708 285326
rect 145656 285262 145708 285268
rect 145668 279970 145696 285262
rect 144656 279942 144716 279970
rect 145024 279942 145084 279970
rect 145452 279942 145696 279970
rect 145760 279970 145788 327655
rect 146116 286544 146168 286550
rect 146116 286486 146168 286492
rect 145760 279942 145820 279970
rect 146128 279834 146156 286486
rect 146496 279970 146524 358090
rect 146864 279970 146892 358158
rect 147496 282328 147548 282334
rect 147496 282270 147548 282276
rect 147508 279970 147536 282270
rect 146496 279942 146556 279970
rect 146864 279942 146924 279970
rect 147292 279942 147536 279970
rect 147600 279970 147628 358226
rect 154948 348492 155000 348498
rect 154948 348434 155000 348440
rect 148324 345092 148376 345098
rect 148324 345034 148376 345040
rect 148336 287910 148364 345034
rect 150900 341624 150952 341630
rect 150900 341566 150952 341572
rect 149428 313948 149480 313954
rect 149428 313890 149480 313896
rect 148324 287904 148376 287910
rect 148324 287846 148376 287852
rect 149060 285048 149112 285054
rect 149060 284990 149112 284996
rect 148968 282464 149020 282470
rect 148968 282406 149020 282412
rect 148232 282396 148284 282402
rect 148232 282338 148284 282344
rect 148244 279970 148272 282338
rect 148598 282160 148654 282169
rect 148598 282095 148654 282104
rect 148612 279970 148640 282095
rect 148980 279970 149008 282406
rect 147600 279942 147660 279970
rect 148028 279942 148272 279970
rect 148396 279942 148640 279970
rect 148764 279942 149008 279970
rect 149072 279970 149100 284990
rect 149440 279970 149468 313890
rect 150532 311160 150584 311166
rect 150532 311102 150584 311108
rect 149796 301504 149848 301510
rect 149796 301446 149848 301452
rect 149808 279970 149836 301446
rect 149980 284980 150032 284986
rect 149980 284922 150032 284928
rect 149992 279970 150020 284922
rect 150544 279970 150572 311102
rect 150912 279970 150940 341566
rect 154580 336048 154632 336054
rect 154580 335990 154632 335996
rect 152372 333328 152424 333334
rect 152372 333270 152424 333276
rect 151268 331900 151320 331906
rect 151268 331842 151320 331848
rect 151280 279970 151308 331842
rect 151636 302932 151688 302938
rect 151636 302874 151688 302880
rect 151648 279970 151676 302874
rect 152004 298784 152056 298790
rect 152004 298726 152056 298732
rect 152016 279970 152044 298726
rect 152384 279970 152412 333270
rect 153844 329112 153896 329118
rect 153844 329054 153896 329060
rect 152740 323672 152792 323678
rect 152740 323614 152792 323620
rect 152752 279970 152780 323614
rect 153108 308508 153160 308514
rect 153108 308450 153160 308456
rect 153120 279970 153148 308450
rect 153476 307080 153528 307086
rect 153476 307022 153528 307028
rect 153488 279970 153516 307022
rect 153856 279970 153884 329054
rect 154212 289196 154264 289202
rect 154212 289138 154264 289144
rect 154224 279970 154252 289138
rect 154592 279970 154620 335990
rect 154960 279970 154988 348434
rect 157616 340332 157668 340338
rect 157616 340274 157668 340280
rect 156420 330608 156472 330614
rect 156420 330550 156472 330556
rect 156052 327820 156104 327826
rect 156052 327762 156104 327768
rect 155684 318096 155736 318102
rect 155684 318038 155736 318044
rect 155316 309800 155368 309806
rect 155316 309742 155368 309748
rect 155328 279970 155356 309742
rect 155696 279970 155724 318038
rect 156064 279970 156092 327762
rect 156236 281852 156288 281858
rect 156236 281794 156288 281800
rect 156248 281654 156276 281794
rect 156236 281648 156288 281654
rect 156236 281590 156288 281596
rect 156432 279970 156460 330550
rect 157156 287904 157208 287910
rect 157156 287846 157208 287852
rect 156788 287700 156840 287706
rect 156788 287642 156840 287648
rect 156800 279970 156828 287642
rect 157168 279970 157196 287846
rect 157628 280242 157656 340274
rect 158260 290488 158312 290494
rect 158260 290430 158312 290436
rect 157892 287768 157944 287774
rect 157892 287710 157944 287716
rect 157582 280214 157656 280242
rect 149072 279942 149132 279970
rect 149440 279942 149500 279970
rect 149808 279942 149868 279970
rect 149992 279942 150236 279970
rect 150544 279942 150604 279970
rect 150912 279942 150972 279970
rect 151280 279942 151340 279970
rect 151648 279942 151708 279970
rect 152016 279942 152076 279970
rect 152384 279942 152444 279970
rect 152752 279942 152812 279970
rect 153120 279942 153180 279970
rect 153488 279942 153548 279970
rect 153856 279942 153916 279970
rect 154224 279942 154284 279970
rect 154592 279942 154652 279970
rect 154960 279942 155020 279970
rect 155328 279942 155388 279970
rect 155696 279942 155756 279970
rect 156064 279942 156124 279970
rect 156432 279942 156492 279970
rect 156800 279942 156860 279970
rect 157168 279942 157228 279970
rect 157582 279956 157610 280214
rect 157904 279970 157932 287710
rect 158272 279970 158300 290430
rect 158628 289264 158680 289270
rect 158628 289206 158680 289212
rect 158640 279970 158668 289206
rect 172980 287564 173032 287570
rect 172980 287506 173032 287512
rect 167092 287496 167144 287502
rect 167092 287438 167144 287444
rect 166908 286476 166960 286482
rect 166908 286418 166960 286424
rect 161020 283484 161072 283490
rect 161020 283426 161072 283432
rect 160100 283416 160152 283422
rect 160100 283358 160152 283364
rect 158904 281988 158956 281994
rect 158904 281930 158956 281936
rect 158812 281920 158864 281926
rect 158812 281862 158864 281868
rect 157904 279942 157964 279970
rect 158272 279942 158332 279970
rect 158640 279942 158700 279970
rect 146128 279806 146188 279834
rect 158824 279614 158852 281862
rect 158916 279970 158944 281930
rect 159180 281852 159232 281858
rect 159180 281794 159232 281800
rect 159192 279970 159220 281794
rect 159548 280492 159600 280498
rect 159548 280434 159600 280440
rect 159560 279970 159588 280434
rect 160112 279970 160140 283358
rect 160284 281648 160336 281654
rect 160284 281590 160336 281596
rect 160296 279970 160324 281590
rect 160652 281580 160704 281586
rect 160652 281522 160704 281528
rect 160664 279970 160692 281522
rect 161032 279970 161060 283426
rect 166264 282600 166316 282606
rect 166264 282542 166316 282548
rect 162860 282532 162912 282538
rect 162860 282474 162912 282480
rect 162124 281784 162176 281790
rect 162124 281726 162176 281732
rect 161572 280356 161624 280362
rect 161572 280298 161624 280304
rect 161584 279970 161612 280298
rect 161756 280288 161808 280294
rect 161756 280230 161808 280236
rect 161768 279970 161796 280230
rect 162136 279970 162164 281726
rect 162492 280832 162544 280838
rect 162492 280774 162544 280780
rect 162504 279970 162532 280774
rect 162872 279970 162900 282474
rect 165068 282124 165120 282130
rect 165068 282066 165120 282072
rect 163964 282056 164016 282062
rect 163964 281998 164016 282004
rect 163596 280424 163648 280430
rect 163596 280366 163648 280372
rect 163458 280220 163510 280226
rect 163458 280162 163510 280168
rect 158916 279942 159068 279970
rect 159192 279942 159436 279970
rect 159560 279942 159804 279970
rect 160112 279942 160172 279970
rect 160296 279942 160540 279970
rect 160664 279942 160908 279970
rect 161032 279942 161276 279970
rect 161584 279942 161644 279970
rect 161768 279942 162012 279970
rect 162136 279942 162380 279970
rect 162504 279942 162748 279970
rect 162872 279942 163116 279970
rect 163470 279956 163498 280162
rect 163608 279970 163636 280366
rect 163976 279970 164004 281998
rect 164332 281920 164384 281926
rect 164332 281862 164384 281868
rect 164344 279970 164372 281862
rect 164700 281716 164752 281722
rect 164700 281658 164752 281664
rect 164712 279970 164740 281658
rect 165080 279970 165108 282066
rect 165666 280220 165718 280226
rect 165666 280162 165718 280168
rect 163608 279942 163852 279970
rect 163976 279942 164220 279970
rect 164344 279942 164588 279970
rect 164712 279942 164956 279970
rect 165080 279942 165324 279970
rect 165678 279956 165706 280162
rect 166276 279970 166304 282542
rect 166632 281580 166684 281586
rect 166632 281522 166684 281528
rect 166644 279970 166672 281522
rect 166920 279970 166948 286418
rect 166060 279942 166304 279970
rect 166428 279942 166672 279970
rect 166796 279942 166948 279970
rect 167104 279970 167132 287438
rect 172612 287428 172664 287434
rect 172612 287370 172664 287376
rect 168840 286408 168892 286414
rect 168840 286350 168892 286356
rect 167736 281716 167788 281722
rect 167736 281658 167788 281664
rect 167748 279970 167776 281658
rect 168104 281648 168156 281654
rect 168104 281590 168156 281596
rect 168116 279970 168144 281590
rect 168196 280628 168248 280634
rect 168196 280570 168248 280576
rect 167104 279942 167164 279970
rect 167532 279942 167776 279970
rect 167900 279942 168144 279970
rect 168208 279834 168236 280570
rect 168852 279970 168880 286350
rect 170680 286340 170732 286346
rect 170680 286282 170732 286288
rect 170312 285116 170364 285122
rect 170312 285058 170364 285064
rect 169668 284436 169720 284442
rect 169668 284378 169720 284384
rect 169576 282056 169628 282062
rect 169576 281998 169628 282004
rect 169208 281852 169260 281858
rect 169208 281794 169260 281800
rect 169220 279970 169248 281794
rect 169588 279970 169616 281998
rect 168636 279942 168880 279970
rect 169004 279942 169248 279970
rect 169372 279942 169616 279970
rect 169680 279970 169708 284378
rect 169760 283552 169812 283558
rect 169760 283494 169812 283500
rect 169772 281654 169800 283494
rect 169760 281648 169812 281654
rect 169760 281590 169812 281596
rect 170324 279970 170352 285058
rect 170692 279970 170720 286282
rect 172428 286272 172480 286278
rect 172428 286214 172480 286220
rect 172152 285048 172204 285054
rect 172152 284990 172204 284996
rect 171416 281988 171468 281994
rect 171416 281930 171468 281936
rect 170956 281920 171008 281926
rect 170956 281862 171008 281868
rect 170968 279970 170996 281862
rect 171428 279970 171456 281930
rect 171784 280424 171836 280430
rect 171784 280366 171836 280372
rect 171796 279970 171824 280366
rect 172164 279970 172192 284990
rect 172440 279970 172468 286214
rect 169680 279942 169740 279970
rect 170108 279942 170352 279970
rect 170476 279942 170720 279970
rect 170844 279942 170996 279970
rect 171212 279942 171456 279970
rect 171580 279942 171824 279970
rect 171948 279942 172192 279970
rect 172316 279942 172468 279970
rect 172624 279970 172652 287370
rect 172992 279970 173020 287506
rect 174360 286204 174412 286210
rect 174360 286146 174412 286152
rect 173808 283416 173860 283422
rect 173808 283358 173860 283364
rect 173716 282532 173768 282538
rect 173716 282474 173768 282480
rect 173624 280492 173676 280498
rect 173624 280434 173676 280440
rect 173636 279970 173664 280434
rect 172624 279942 172684 279970
rect 172992 279942 173052 279970
rect 173420 279942 173664 279970
rect 173728 279970 173756 282474
rect 173820 282266 173848 283358
rect 173808 282260 173860 282266
rect 173808 282202 173860 282208
rect 174372 279970 174400 286146
rect 176200 286136 176252 286142
rect 176200 286078 176252 286084
rect 175832 284980 175884 284986
rect 175832 284922 175884 284928
rect 174912 283484 174964 283490
rect 174912 283426 174964 283432
rect 174924 282198 174952 283426
rect 174912 282192 174964 282198
rect 174912 282134 174964 282140
rect 175004 282124 175056 282130
rect 175004 282066 175056 282072
rect 174728 281784 174780 281790
rect 174728 281726 174780 281732
rect 174740 279970 174768 281726
rect 175016 279970 175044 282066
rect 175186 281888 175242 281897
rect 175186 281823 175242 281832
rect 175096 280832 175148 280838
rect 175200 280809 175228 281823
rect 175096 280774 175148 280780
rect 175186 280800 175242 280809
rect 173728 279942 173788 279970
rect 174156 279942 174400 279970
rect 174524 279942 174768 279970
rect 174892 279942 175044 279970
rect 175108 279970 175136 280774
rect 175186 280735 175242 280744
rect 175844 279970 175872 284922
rect 175922 281752 175978 281761
rect 175922 281687 175978 281696
rect 175936 280945 175964 281687
rect 175922 280936 175978 280945
rect 175922 280871 175978 280880
rect 176212 279970 176240 286078
rect 176672 282470 176700 700266
rect 177210 597000 177266 597009
rect 177210 596935 177266 596944
rect 177224 296070 177252 596935
rect 177212 296064 177264 296070
rect 177212 296006 177264 296012
rect 176752 287632 176804 287638
rect 176752 287574 176804 287580
rect 176660 282464 176712 282470
rect 176660 282406 176712 282412
rect 176568 281648 176620 281654
rect 176568 281590 176620 281596
rect 176580 279970 176608 281590
rect 176764 280242 176792 287574
rect 177316 285258 177344 700266
rect 177408 285326 177436 700402
rect 177948 597032 178000 597038
rect 177948 596974 178000 596980
rect 177856 596692 177908 596698
rect 177856 596634 177908 596640
rect 177764 596488 177816 596494
rect 177764 596430 177816 596436
rect 177580 596420 177632 596426
rect 177580 596362 177632 596368
rect 177488 596284 177540 596290
rect 177488 596226 177540 596232
rect 177500 290873 177528 596226
rect 177592 292058 177620 596362
rect 177672 596352 177724 596358
rect 177672 596294 177724 596300
rect 177580 292052 177632 292058
rect 177580 291994 177632 292000
rect 177486 290864 177542 290873
rect 177486 290799 177542 290808
rect 177684 290737 177712 596294
rect 177776 293622 177804 596430
rect 177868 295118 177896 596634
rect 177960 296274 177988 596974
rect 177948 296268 178000 296274
rect 177948 296210 178000 296216
rect 177856 295112 177908 295118
rect 177856 295054 177908 295060
rect 177764 293616 177816 293622
rect 177764 293558 177816 293564
rect 177670 290728 177726 290737
rect 177670 290663 177726 290672
rect 177396 285320 177448 285326
rect 177396 285262 177448 285268
rect 177304 285252 177356 285258
rect 177304 285194 177356 285200
rect 178052 282690 178080 700538
rect 178224 700528 178276 700534
rect 178224 700470 178276 700476
rect 178132 700392 178184 700398
rect 178132 700334 178184 700340
rect 178144 282849 178172 700334
rect 178130 282840 178186 282849
rect 178130 282775 178186 282784
rect 178052 282662 178172 282690
rect 178040 282600 178092 282606
rect 178040 282542 178092 282548
rect 177948 282464 178000 282470
rect 177948 282406 178000 282412
rect 177304 280356 177356 280362
rect 177304 280298 177356 280304
rect 175108 279942 175260 279970
rect 175628 279942 175872 279970
rect 175996 279942 176240 279970
rect 176364 279942 176608 279970
rect 176718 280214 176792 280242
rect 176718 279956 176746 280214
rect 177316 279970 177344 280298
rect 177960 279970 177988 282406
rect 178052 280974 178080 282542
rect 178144 282334 178172 282662
rect 178236 282402 178264 700470
rect 178328 358222 178356 700674
rect 178408 700664 178460 700670
rect 178408 700606 178460 700612
rect 178420 358290 178448 700606
rect 186964 700392 187016 700398
rect 186964 700334 187016 700340
rect 178498 679144 178554 679153
rect 178498 679079 178554 679088
rect 178512 560289 178540 679079
rect 178960 597100 179012 597106
rect 178960 597042 179012 597048
rect 178776 596964 178828 596970
rect 178776 596906 178828 596912
rect 178684 596760 178736 596766
rect 178684 596702 178736 596708
rect 178498 560280 178554 560289
rect 178498 560215 178554 560224
rect 178500 444372 178552 444378
rect 178500 444314 178552 444320
rect 178512 443290 178540 444314
rect 178500 443284 178552 443290
rect 178500 443226 178552 443232
rect 178512 439249 178540 443226
rect 178498 439240 178554 439249
rect 178498 439175 178554 439184
rect 178408 358284 178460 358290
rect 178408 358226 178460 358232
rect 178316 358216 178368 358222
rect 178316 358158 178368 358164
rect 178696 294982 178724 596702
rect 178684 294976 178736 294982
rect 178684 294918 178736 294924
rect 178788 294778 178816 596906
rect 178868 596828 178920 596834
rect 178868 596770 178920 596776
rect 178880 294914 178908 596770
rect 178972 296206 179000 597042
rect 182824 596896 182876 596902
rect 182824 596838 182876 596844
rect 180064 596556 180116 596562
rect 180064 596498 180116 596504
rect 179050 560280 179106 560289
rect 179050 560215 179106 560224
rect 179064 559201 179092 560215
rect 179050 559192 179106 559201
rect 179050 559127 179106 559136
rect 179064 453354 179092 559127
rect 179052 453348 179104 453354
rect 179052 453290 179104 453296
rect 179064 444378 179092 453290
rect 179052 444372 179104 444378
rect 179052 444314 179104 444320
rect 178960 296200 179012 296206
rect 178960 296142 179012 296148
rect 178868 294908 178920 294914
rect 178868 294850 178920 294856
rect 178776 294772 178828 294778
rect 178776 294714 178828 294720
rect 180076 291990 180104 596498
rect 180154 487248 180210 487257
rect 180154 487183 180210 487192
rect 180168 447098 180196 487183
rect 180156 447092 180208 447098
rect 180156 447034 180208 447040
rect 182836 294846 182864 596838
rect 182916 470620 182968 470626
rect 182916 470562 182968 470568
rect 182824 294840 182876 294846
rect 182824 294782 182876 294788
rect 182928 292126 182956 470562
rect 186976 358154 187004 700334
rect 192484 696992 192536 696998
rect 192484 696934 192536 696940
rect 191104 596624 191156 596630
rect 191104 596566 191156 596572
rect 188344 590708 188396 590714
rect 188344 590650 188396 590656
rect 186964 358148 187016 358154
rect 186964 358090 187016 358096
rect 188356 305658 188384 590650
rect 188436 456816 188488 456822
rect 188436 456758 188488 456764
rect 188344 305652 188396 305658
rect 188344 305594 188396 305600
rect 182916 292120 182968 292126
rect 182916 292062 182968 292068
rect 180064 291984 180116 291990
rect 180064 291926 180116 291932
rect 182916 287360 182968 287366
rect 181810 287328 181866 287337
rect 182916 287302 182968 287308
rect 181810 287263 181866 287272
rect 181352 286068 181404 286074
rect 181352 286010 181404 286016
rect 179236 284912 179288 284918
rect 179236 284854 179288 284860
rect 179144 284368 179196 284374
rect 179144 284310 179196 284316
rect 178316 283756 178368 283762
rect 178316 283698 178368 283704
rect 178328 282538 178356 283698
rect 178316 282532 178368 282538
rect 178316 282474 178368 282480
rect 178224 282396 178276 282402
rect 178224 282338 178276 282344
rect 178132 282328 178184 282334
rect 178132 282270 178184 282276
rect 178408 282192 178460 282198
rect 178408 282134 178460 282140
rect 178040 280968 178092 280974
rect 178040 280910 178092 280916
rect 178420 279970 178448 282134
rect 178774 281752 178830 281761
rect 178774 281687 178830 281696
rect 178788 279970 178816 281687
rect 179156 279970 179184 284310
rect 177100 279942 177344 279970
rect 177836 279942 177988 279970
rect 178204 279942 178448 279970
rect 178572 279942 178816 279970
rect 178940 279942 179184 279970
rect 179248 279834 179276 284854
rect 179880 284844 179932 284850
rect 179880 284786 179932 284792
rect 179420 281580 179472 281586
rect 179420 281522 179472 281528
rect 168208 279806 168268 279834
rect 179248 279806 179308 279834
rect 179432 279818 179460 281522
rect 179892 279970 179920 284786
rect 180248 282396 180300 282402
rect 180248 282338 180300 282344
rect 180260 279970 180288 282338
rect 180708 280560 180760 280566
rect 180708 280502 180760 280508
rect 179676 279942 179920 279970
rect 180044 279942 180288 279970
rect 180720 279970 180748 280502
rect 181364 279970 181392 286010
rect 181720 282260 181772 282266
rect 181720 282202 181772 282208
rect 181732 279970 181760 282202
rect 180720 279942 180780 279970
rect 181148 279942 181392 279970
rect 181516 279942 181760 279970
rect 181824 279970 181852 287263
rect 182456 286000 182508 286006
rect 182456 285942 182508 285948
rect 182468 279970 182496 285942
rect 182824 285932 182876 285938
rect 182824 285874 182876 285880
rect 182836 279970 182864 285874
rect 181824 279942 181884 279970
rect 182252 279942 182496 279970
rect 182620 279942 182864 279970
rect 182928 279970 182956 287302
rect 184388 287292 184440 287298
rect 184388 287234 184440 287240
rect 184296 285864 184348 285870
rect 184296 285806 184348 285812
rect 183466 282160 183522 282169
rect 183466 282095 183522 282104
rect 183480 279970 183508 282095
rect 184308 279970 184336 285806
rect 182928 279942 182988 279970
rect 183356 279942 183508 279970
rect 184092 279942 184336 279970
rect 184400 279970 184428 287234
rect 187332 287224 187384 287230
rect 187332 287166 187384 287172
rect 187698 287192 187754 287201
rect 185768 285796 185820 285802
rect 185768 285738 185820 285744
rect 185400 284776 185452 284782
rect 185400 284718 185452 284724
rect 184756 281104 184808 281110
rect 184756 281046 184808 281052
rect 184768 279970 184796 281046
rect 185412 279970 185440 284718
rect 185582 281616 185638 281625
rect 185582 281551 185638 281560
rect 185596 280838 185624 281551
rect 185492 280832 185544 280838
rect 185492 280774 185544 280780
rect 185584 280832 185636 280838
rect 185584 280774 185636 280780
rect 185504 280362 185532 280774
rect 185492 280356 185544 280362
rect 185492 280298 185544 280304
rect 185780 279970 185808 285738
rect 187240 285728 187292 285734
rect 187240 285670 187292 285676
rect 186872 284708 186924 284714
rect 186872 284650 186924 284656
rect 186136 282328 186188 282334
rect 186136 282270 186188 282276
rect 186148 279970 186176 282270
rect 186226 281616 186282 281625
rect 186226 281551 186282 281560
rect 184400 279942 184460 279970
rect 184768 279942 184828 279970
rect 185196 279942 185440 279970
rect 185564 279942 185808 279970
rect 185932 279942 186176 279970
rect 186240 279970 186268 281551
rect 186884 279970 186912 284650
rect 187252 279970 187280 285670
rect 186240 279942 186300 279970
rect 186668 279942 186912 279970
rect 187036 279942 187280 279970
rect 187344 279970 187372 287166
rect 187698 287127 187754 287136
rect 187712 279970 187740 287127
rect 188448 285190 188476 456758
rect 191116 295050 191144 596566
rect 192116 356244 192168 356250
rect 192116 356186 192168 356192
rect 191196 351960 191248 351966
rect 191196 351902 191248 351908
rect 191104 295044 191156 295050
rect 191104 294986 191156 294992
rect 191208 287842 191236 351902
rect 191380 351212 191432 351218
rect 191380 351154 191432 351160
rect 191196 287836 191248 287842
rect 191196 287778 191248 287784
rect 189906 287464 189962 287473
rect 189906 287399 189962 287408
rect 189540 287156 189592 287162
rect 189540 287098 189592 287104
rect 188436 285184 188488 285190
rect 188436 285126 188488 285132
rect 188344 284640 188396 284646
rect 188344 284582 188396 284588
rect 187792 283688 187844 283694
rect 187792 283630 187844 283636
rect 187804 282470 187832 283630
rect 187792 282464 187844 282470
rect 187792 282406 187844 282412
rect 187884 282396 187936 282402
rect 187884 282338 187936 282344
rect 187344 279942 187404 279970
rect 187712 279942 187772 279970
rect 179420 279812 179472 279818
rect 179420 279754 179472 279760
rect 187896 279750 187924 282338
rect 188356 279970 188384 284582
rect 189448 284572 189500 284578
rect 189448 284514 189500 284520
rect 188986 282024 189042 282033
rect 188986 281959 189042 281968
rect 188712 281580 188764 281586
rect 188712 281522 188764 281528
rect 188724 279970 188752 281522
rect 189000 279970 189028 281959
rect 189460 279970 189488 284514
rect 188140 279942 188384 279970
rect 188508 279942 188752 279970
rect 188876 279942 189028 279970
rect 189244 279942 189488 279970
rect 189552 279970 189580 287098
rect 189920 279970 189948 287399
rect 190644 287088 190696 287094
rect 190644 287030 190696 287036
rect 190276 284504 190328 284510
rect 190276 284446 190328 284452
rect 190288 279970 190316 284446
rect 190656 279970 190684 287030
rect 191286 281888 191342 281897
rect 191286 281823 191342 281832
rect 191300 279970 191328 281823
rect 189552 279942 189612 279970
rect 189920 279942 189980 279970
rect 190288 279942 190348 279970
rect 190656 279942 190716 279970
rect 191084 279942 191328 279970
rect 191392 279970 191420 351154
rect 192024 326460 192076 326466
rect 192024 326402 192076 326408
rect 191748 291848 191800 291854
rect 191748 291790 191800 291796
rect 191656 282328 191708 282334
rect 191656 282270 191708 282276
rect 191668 280906 191696 282270
rect 191656 280900 191708 280906
rect 191656 280842 191708 280848
rect 191760 279970 191788 291790
rect 192036 282878 192064 326402
rect 192024 282872 192076 282878
rect 192024 282814 192076 282820
rect 192128 279970 192156 356186
rect 192496 318238 192524 696934
rect 192576 685908 192628 685914
rect 192576 685850 192628 685856
rect 192588 607918 192616 685850
rect 192576 607912 192628 607918
rect 192576 607854 192628 607860
rect 200764 596216 200816 596222
rect 200764 596158 200816 596164
rect 193864 576904 193916 576910
rect 193864 576846 193916 576852
rect 192852 330676 192904 330682
rect 192852 330618 192904 330624
rect 192484 318232 192536 318238
rect 192484 318174 192536 318180
rect 192300 282872 192352 282878
rect 192300 282814 192352 282820
rect 192312 279970 192340 282814
rect 192864 279970 192892 330618
rect 193876 323746 193904 576846
rect 200120 358080 200172 358086
rect 200120 358022 200172 358028
rect 196532 356312 196584 356318
rect 196532 356254 196584 356260
rect 195428 337408 195480 337414
rect 195428 337350 195480 337356
rect 193864 323740 193916 323746
rect 193864 323682 193916 323688
rect 194324 322312 194376 322318
rect 194324 322254 194376 322260
rect 193956 312588 194008 312594
rect 193956 312530 194008 312536
rect 193588 298852 193640 298858
rect 193588 298794 193640 298800
rect 193220 294636 193272 294642
rect 193220 294578 193272 294584
rect 193232 279970 193260 294578
rect 193600 279970 193628 298794
rect 193968 279970 193996 312530
rect 194336 279970 194364 322254
rect 195060 308440 195112 308446
rect 195060 308382 195112 308388
rect 194692 295996 194744 296002
rect 194692 295938 194744 295944
rect 194704 279970 194732 295938
rect 195072 279970 195100 308382
rect 195440 279970 195468 337350
rect 195796 323604 195848 323610
rect 195796 323546 195848 323552
rect 195808 279970 195836 323546
rect 196164 297424 196216 297430
rect 196164 297366 196216 297372
rect 196176 279970 196204 297366
rect 196544 279970 196572 356254
rect 198372 356108 198424 356114
rect 198372 356050 198424 356056
rect 197636 352572 197688 352578
rect 197636 352514 197688 352520
rect 196900 316736 196952 316742
rect 196900 316678 196952 316684
rect 196912 279970 196940 316678
rect 197268 294704 197320 294710
rect 197268 294646 197320 294652
rect 197280 279970 197308 294646
rect 197648 279970 197676 352514
rect 198004 311228 198056 311234
rect 198004 311170 198056 311176
rect 198016 279970 198044 311170
rect 198384 279970 198412 356050
rect 199844 355360 199896 355366
rect 199844 355302 199896 355308
rect 198740 354000 198792 354006
rect 198740 353942 198792 353948
rect 198752 279970 198780 353942
rect 199476 327888 199528 327894
rect 199476 327830 199528 327836
rect 199108 309868 199160 309874
rect 199108 309810 199160 309816
rect 199120 279970 199148 309810
rect 199488 279970 199516 327830
rect 199856 279970 199884 355302
rect 200132 282878 200160 358022
rect 200580 329180 200632 329186
rect 200580 329122 200632 329128
rect 200212 291916 200264 291922
rect 200212 291858 200264 291864
rect 200120 282872 200172 282878
rect 200120 282814 200172 282820
rect 200224 279970 200252 291858
rect 200592 279970 200620 329122
rect 200776 293282 200804 596158
rect 200948 565480 201000 565486
rect 200948 565422 201000 565428
rect 200856 565412 200908 565418
rect 200856 565354 200908 565360
rect 200868 293758 200896 565354
rect 200856 293752 200908 293758
rect 200856 293694 200908 293700
rect 200960 293690 200988 565422
rect 201040 565344 201092 565350
rect 201040 565286 201092 565292
rect 201052 293894 201080 565286
rect 201040 293888 201092 293894
rect 201040 293830 201092 293836
rect 200948 293684 201000 293690
rect 200948 293626 201000 293632
rect 201316 293344 201368 293350
rect 201316 293286 201368 293292
rect 200764 293276 200816 293282
rect 200764 293218 200816 293224
rect 200764 282872 200816 282878
rect 200764 282814 200816 282820
rect 200776 279970 200804 282814
rect 201328 279970 201356 293286
rect 201512 286550 201540 702986
rect 218992 700398 219020 703520
rect 235184 700777 235212 703520
rect 235170 700768 235226 700777
rect 235170 700703 235226 700712
rect 267660 700641 267688 703520
rect 267646 700632 267702 700641
rect 267646 700567 267702 700576
rect 283852 700466 283880 703520
rect 300136 700505 300164 703520
rect 300122 700496 300178 700505
rect 283840 700460 283892 700466
rect 300122 700431 300178 700440
rect 283840 700402 283892 700408
rect 218980 700392 219032 700398
rect 332520 700369 332548 703520
rect 218980 700334 219032 700340
rect 332506 700360 332562 700369
rect 348804 700330 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 360844 700392 360896 700398
rect 360844 700334 360896 700340
rect 332506 700295 332562 700304
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 350998 685944 351054 685953
rect 350998 685879 351000 685888
rect 351052 685879 351054 685888
rect 351000 685850 351052 685856
rect 358818 679008 358874 679017
rect 358818 678943 358874 678952
rect 217230 636848 217286 636857
rect 217230 636783 217286 636792
rect 217138 635896 217194 635905
rect 217138 635831 217194 635840
rect 216678 608288 216734 608297
rect 216678 608223 216734 608232
rect 213920 607912 213972 607918
rect 213920 607854 213972 607860
rect 213932 607374 213960 607854
rect 216692 607374 216720 608223
rect 213920 607368 213972 607374
rect 213920 607310 213972 607316
rect 216680 607368 216732 607374
rect 216680 607310 216732 607316
rect 213550 597408 213606 597417
rect 213550 597343 213606 597352
rect 211066 597000 211122 597009
rect 211066 596935 211122 596944
rect 210976 594244 211028 594250
rect 210976 594186 211028 594192
rect 204076 565752 204128 565758
rect 204076 565694 204128 565700
rect 203892 565684 203944 565690
rect 203892 565626 203944 565632
rect 203800 565616 203852 565622
rect 203800 565558 203852 565564
rect 203708 565548 203760 565554
rect 203708 565490 203760 565496
rect 203616 565208 203668 565214
rect 203616 565150 203668 565156
rect 203524 565140 203576 565146
rect 203524 565082 203576 565088
rect 203156 356176 203208 356182
rect 203156 356118 203208 356124
rect 202972 349852 203024 349858
rect 202972 349794 203024 349800
rect 202420 344412 202472 344418
rect 202420 344354 202472 344360
rect 202052 314016 202104 314022
rect 202052 313958 202104 313964
rect 201868 296132 201920 296138
rect 201868 296074 201920 296080
rect 201500 286544 201552 286550
rect 201500 286486 201552 286492
rect 201880 279970 201908 296074
rect 191392 279942 191452 279970
rect 191760 279942 191820 279970
rect 192128 279942 192188 279970
rect 192312 279942 192556 279970
rect 192864 279942 192924 279970
rect 193232 279942 193292 279970
rect 193600 279942 193660 279970
rect 193968 279942 194028 279970
rect 194336 279942 194396 279970
rect 194704 279942 194764 279970
rect 195072 279942 195132 279970
rect 195440 279942 195500 279970
rect 195808 279942 195868 279970
rect 196176 279942 196236 279970
rect 196544 279942 196604 279970
rect 196912 279942 196972 279970
rect 197280 279942 197340 279970
rect 197648 279942 197708 279970
rect 198016 279942 198076 279970
rect 198384 279942 198444 279970
rect 198752 279942 198812 279970
rect 199120 279942 199180 279970
rect 199488 279942 199548 279970
rect 199856 279942 199916 279970
rect 200224 279942 200284 279970
rect 200592 279942 200652 279970
rect 200776 279942 201020 279970
rect 201328 279942 201388 279970
rect 201756 279942 201908 279970
rect 202064 279970 202092 313958
rect 202432 279970 202460 344354
rect 202788 315376 202840 315382
rect 202788 315318 202840 315324
rect 202800 279970 202828 315318
rect 202984 282878 203012 349794
rect 203064 318164 203116 318170
rect 203064 318106 203116 318112
rect 202972 282872 203024 282878
rect 202972 282814 203024 282820
rect 203076 282810 203104 318106
rect 203064 282804 203116 282810
rect 203064 282746 203116 282752
rect 203168 279970 203196 356118
rect 203536 285258 203564 565082
rect 203628 291009 203656 565150
rect 203720 293554 203748 565490
rect 203708 293548 203760 293554
rect 203708 293490 203760 293496
rect 203812 293486 203840 565558
rect 203800 293480 203852 293486
rect 203800 293422 203852 293428
rect 203904 293418 203932 565626
rect 203984 565276 204036 565282
rect 203984 565218 204036 565224
rect 203996 293962 204024 565218
rect 203984 293956 204036 293962
rect 203984 293898 204036 293904
rect 203892 293412 203944 293418
rect 203892 293354 203944 293360
rect 204088 293350 204116 565694
rect 210698 477456 210754 477465
rect 210698 477391 210754 477400
rect 210422 477320 210478 477329
rect 210422 477255 210478 477264
rect 207020 477216 207072 477222
rect 207020 477158 207072 477164
rect 208308 477216 208360 477222
rect 208308 477158 208360 477164
rect 207032 476406 207060 477158
rect 207020 476400 207072 476406
rect 207020 476342 207072 476348
rect 206560 448180 206612 448186
rect 206560 448122 206612 448128
rect 206468 447976 206520 447982
rect 206468 447918 206520 447924
rect 206376 447908 206428 447914
rect 206376 447850 206428 447856
rect 206284 447840 206336 447846
rect 206284 447782 206336 447788
rect 205364 348560 205416 348566
rect 205364 348502 205416 348508
rect 204628 340264 204680 340270
rect 204628 340206 204680 340212
rect 204260 300144 204312 300150
rect 204260 300086 204312 300092
rect 204076 293344 204128 293350
rect 204076 293286 204128 293292
rect 203614 291000 203670 291009
rect 203614 290935 203670 290944
rect 203524 285252 203576 285258
rect 203524 285194 203576 285200
rect 203340 282872 203392 282878
rect 203340 282814 203392 282820
rect 203352 279970 203380 282814
rect 203708 282804 203760 282810
rect 203708 282746 203760 282752
rect 203720 279970 203748 282746
rect 204272 279970 204300 300086
rect 204640 279970 204668 340206
rect 204996 301572 205048 301578
rect 204996 301514 205048 301520
rect 205008 279970 205036 301514
rect 205376 279970 205404 348502
rect 206100 347132 206152 347138
rect 206100 347074 206152 347080
rect 206008 304292 206060 304298
rect 206008 304234 206060 304240
rect 205732 303000 205784 303006
rect 205732 302942 205784 302948
rect 205744 279970 205772 302942
rect 206020 282878 206048 304234
rect 206008 282872 206060 282878
rect 206008 282814 206060 282820
rect 206112 279970 206140 347074
rect 206296 284730 206324 447782
rect 206388 285190 206416 447850
rect 206480 287910 206508 447918
rect 206572 290426 206600 448122
rect 206652 448112 206704 448118
rect 206652 448054 206704 448060
rect 206560 290420 206612 290426
rect 206560 290362 206612 290368
rect 206664 290358 206692 448054
rect 206744 448044 206796 448050
rect 206744 447986 206796 447992
rect 206652 290352 206704 290358
rect 206652 290294 206704 290300
rect 206756 290290 206784 447986
rect 208320 355842 208348 477158
rect 210436 476649 210464 477255
rect 210422 476640 210478 476649
rect 210422 476575 210478 476584
rect 208952 474088 209004 474094
rect 208952 474030 209004 474036
rect 208584 445052 208636 445058
rect 208584 444994 208636 445000
rect 208308 355836 208360 355842
rect 208308 355778 208360 355784
rect 207940 342916 207992 342922
rect 207940 342858 207992 342864
rect 207572 341692 207624 341698
rect 207572 341634 207624 341640
rect 206836 320952 206888 320958
rect 206836 320894 206888 320900
rect 206744 290284 206796 290290
rect 206744 290226 206796 290232
rect 206468 287904 206520 287910
rect 206468 287846 206520 287852
rect 206376 285184 206428 285190
rect 206376 285126 206428 285132
rect 206296 284702 206416 284730
rect 206284 282872 206336 282878
rect 206284 282814 206336 282820
rect 206296 279970 206324 282814
rect 206388 282402 206416 284702
rect 206376 282396 206428 282402
rect 206376 282338 206428 282344
rect 206848 279970 206876 320894
rect 207204 307148 207256 307154
rect 207204 307090 207256 307096
rect 207216 279970 207244 307090
rect 207584 279970 207612 341634
rect 207952 279970 207980 342858
rect 208308 291848 208360 291854
rect 208308 291790 208360 291796
rect 208320 279970 208348 291790
rect 208596 282878 208624 444994
rect 208964 359650 208992 474030
rect 210332 474020 210384 474026
rect 210332 473962 210384 473968
rect 210148 449268 210200 449274
rect 210148 449210 210200 449216
rect 209228 448520 209280 448526
rect 209228 448462 209280 448468
rect 209044 448384 209096 448390
rect 209044 448326 209096 448332
rect 208952 359644 209004 359650
rect 208952 359586 209004 359592
rect 208674 294536 208730 294545
rect 208674 294471 208730 294480
rect 208584 282872 208636 282878
rect 208584 282814 208636 282820
rect 208688 279970 208716 294471
rect 209056 290766 209084 448326
rect 209136 447704 209188 447710
rect 209136 447646 209188 447652
rect 209044 290760 209096 290766
rect 209044 290702 209096 290708
rect 209148 290222 209176 447646
rect 209240 290630 209268 448462
rect 209412 448452 209464 448458
rect 209412 448394 209464 448400
rect 209320 447772 209372 447778
rect 209320 447714 209372 447720
rect 209228 290624 209280 290630
rect 209228 290566 209280 290572
rect 209332 290562 209360 447714
rect 209424 290698 209452 448394
rect 209596 448316 209648 448322
rect 209596 448258 209648 448264
rect 209504 448248 209556 448254
rect 209504 448190 209556 448196
rect 209516 290902 209544 448190
rect 209504 290896 209556 290902
rect 209504 290838 209556 290844
rect 209608 290834 209636 448258
rect 209688 444916 209740 444922
rect 209688 444858 209740 444864
rect 209700 290970 209728 444858
rect 209780 315376 209832 315382
rect 209780 315318 209832 315324
rect 209688 290964 209740 290970
rect 209688 290906 209740 290912
rect 209596 290828 209648 290834
rect 209596 290770 209648 290776
rect 209412 290692 209464 290698
rect 209412 290634 209464 290640
rect 209320 290556 209372 290562
rect 209320 290498 209372 290504
rect 209136 290216 209188 290222
rect 209136 290158 209188 290164
rect 208860 282872 208912 282878
rect 208860 282814 208912 282820
rect 209226 282840 209282 282849
rect 208872 279970 208900 282814
rect 209226 282775 209282 282784
rect 209240 279970 209268 282775
rect 209792 279970 209820 315318
rect 210160 279970 210188 449210
rect 210344 359718 210372 473962
rect 210332 359712 210384 359718
rect 210332 359654 210384 359660
rect 210436 355162 210464 476575
rect 210514 476504 210570 476513
rect 210514 476439 210570 476448
rect 210608 476468 210660 476474
rect 210528 356046 210556 476439
rect 210608 476410 210660 476416
rect 210516 356040 210568 356046
rect 210516 355982 210568 355988
rect 210620 355910 210648 476410
rect 210712 476377 210740 477391
rect 210882 477184 210938 477193
rect 210882 477119 210938 477128
rect 210698 476368 210754 476377
rect 210698 476303 210754 476312
rect 210792 476332 210844 476338
rect 210712 355978 210740 476303
rect 210792 476274 210844 476280
rect 210700 355972 210752 355978
rect 210700 355914 210752 355920
rect 210608 355904 210660 355910
rect 210608 355846 210660 355852
rect 210804 355638 210832 476274
rect 210792 355632 210844 355638
rect 210792 355574 210844 355580
rect 210424 355156 210476 355162
rect 210424 355098 210476 355104
rect 210896 351830 210924 477119
rect 210988 359922 211016 594186
rect 210976 359916 211028 359922
rect 210976 359858 211028 359864
rect 211080 359310 211108 596935
rect 212356 594312 212408 594318
rect 212356 594254 212408 594260
rect 211712 476740 211764 476746
rect 211712 476682 211764 476688
rect 211724 476202 211752 476682
rect 211712 476196 211764 476202
rect 211712 476138 211764 476144
rect 211068 359304 211120 359310
rect 211068 359246 211120 359252
rect 210884 351824 210936 351830
rect 210884 351766 210936 351772
rect 211724 344622 211752 476138
rect 212264 445732 212316 445738
rect 212264 445674 212316 445680
rect 212172 445664 212224 445670
rect 212172 445606 212224 445612
rect 211988 445596 212040 445602
rect 211988 445538 212040 445544
rect 211804 445528 211856 445534
rect 211804 445470 211856 445476
rect 211712 344616 211764 344622
rect 211712 344558 211764 344564
rect 211160 340944 211212 340950
rect 211160 340886 211212 340892
rect 210884 329112 210936 329118
rect 210884 329054 210936 329060
rect 210698 282840 210754 282849
rect 210698 282775 210754 282784
rect 210712 279970 210740 282775
rect 202064 279942 202124 279970
rect 202432 279942 202492 279970
rect 202800 279942 202860 279970
rect 203168 279942 203228 279970
rect 203352 279942 203596 279970
rect 203720 279942 203964 279970
rect 204272 279942 204332 279970
rect 204640 279942 204700 279970
rect 205008 279942 205068 279970
rect 205376 279942 205436 279970
rect 205744 279942 205804 279970
rect 206112 279942 206172 279970
rect 206296 279942 206540 279970
rect 206848 279942 206908 279970
rect 207216 279942 207276 279970
rect 207584 279942 207644 279970
rect 207952 279942 208012 279970
rect 208320 279942 208380 279970
rect 208688 279942 208748 279970
rect 208872 279942 209116 279970
rect 209240 279942 209484 279970
rect 209792 279942 209852 279970
rect 210160 279942 210220 279970
rect 210588 279942 210740 279970
rect 210896 279970 210924 329054
rect 211172 287054 211200 340886
rect 211816 287774 211844 445470
rect 211896 445460 211948 445466
rect 211896 445402 211948 445408
rect 211908 287842 211936 445402
rect 211896 287836 211948 287842
rect 211896 287778 211948 287784
rect 211804 287768 211856 287774
rect 211804 287710 211856 287716
rect 212000 287706 212028 445538
rect 212080 444984 212132 444990
rect 212080 444926 212132 444932
rect 212092 291038 212120 444926
rect 212184 291174 212212 445606
rect 212172 291168 212224 291174
rect 212172 291110 212224 291116
rect 212276 291106 212304 445674
rect 212368 359553 212396 594254
rect 212448 594108 212500 594114
rect 212448 594050 212500 594056
rect 212460 359854 212488 594050
rect 213366 477320 213422 477329
rect 213366 477255 213422 477264
rect 213274 477048 213330 477057
rect 213274 476983 213330 476992
rect 213182 476912 213238 476921
rect 213182 476847 213238 476856
rect 213092 474292 213144 474298
rect 213092 474234 213144 474240
rect 212540 449200 212592 449206
rect 212540 449142 212592 449148
rect 212448 359848 212500 359854
rect 212448 359790 212500 359796
rect 212354 359544 212410 359553
rect 212354 359479 212410 359488
rect 212356 345024 212408 345030
rect 212356 344966 212408 344972
rect 212368 344622 212396 344966
rect 212356 344616 212408 344622
rect 212356 344558 212408 344564
rect 212264 291100 212316 291106
rect 212264 291042 212316 291048
rect 212080 291032 212132 291038
rect 212080 290974 212132 290980
rect 211988 287700 212040 287706
rect 211988 287642 212040 287648
rect 211172 287026 211844 287054
rect 211526 282840 211582 282849
rect 211526 282775 211582 282784
rect 211540 279970 211568 282775
rect 211618 282704 211674 282713
rect 211618 282639 211674 282648
rect 210896 279942 210956 279970
rect 211324 279942 211568 279970
rect 211632 279834 211660 282639
rect 211816 279970 211844 287026
rect 212368 279970 212396 344558
rect 212552 282878 212580 449142
rect 213104 359514 213132 474234
rect 213092 359508 213144 359514
rect 213092 359450 213144 359456
rect 212724 350600 212776 350606
rect 212724 350542 212776 350548
rect 212540 282872 212592 282878
rect 212540 282814 212592 282820
rect 212736 279970 212764 350542
rect 213196 342242 213224 476847
rect 213288 356017 213316 476983
rect 213380 476785 213408 477255
rect 213366 476776 213422 476785
rect 213366 476711 213422 476720
rect 213274 356008 213330 356017
rect 213274 355943 213330 355952
rect 213380 351898 213408 476711
rect 213460 476264 213512 476270
rect 213460 476206 213512 476212
rect 213368 351892 213420 351898
rect 213368 351834 213420 351840
rect 213380 350606 213408 351834
rect 213368 350600 213420 350606
rect 213368 350542 213420 350548
rect 213472 350538 213500 476206
rect 213564 358329 213592 597343
rect 213642 594552 213698 594561
rect 213642 594487 213698 594496
rect 213550 358320 213606 358329
rect 213550 358255 213606 358264
rect 213656 355881 213684 594487
rect 213734 594416 213790 594425
rect 213734 594351 213790 594360
rect 213642 355872 213698 355881
rect 213642 355807 213698 355816
rect 213748 355745 213776 594351
rect 213826 594280 213882 594289
rect 213826 594215 213882 594224
rect 213734 355736 213790 355745
rect 213734 355671 213790 355680
rect 213840 355609 213868 594215
rect 213932 567225 213960 607310
rect 214748 597168 214800 597174
rect 214748 597110 214800 597116
rect 214564 594584 214616 594590
rect 214564 594526 214616 594532
rect 214472 594448 214524 594454
rect 214472 594390 214524 594396
rect 214380 594040 214432 594046
rect 214380 593982 214432 593988
rect 213918 567216 213974 567225
rect 213918 567151 213920 567160
rect 213972 567151 213974 567160
rect 213920 567122 213972 567128
rect 214392 477426 214420 593982
rect 214380 477420 214432 477426
rect 214380 477362 214432 477368
rect 214392 476406 214420 477362
rect 214484 476513 214512 594390
rect 214576 477426 214604 594526
rect 214656 594516 214708 594522
rect 214656 594458 214708 594464
rect 214564 477420 214616 477426
rect 214564 477362 214616 477368
rect 214470 476504 214526 476513
rect 214576 476474 214604 477362
rect 214470 476439 214526 476448
rect 214564 476468 214616 476474
rect 214564 476410 214616 476416
rect 214380 476400 214432 476406
rect 214668 476377 214696 594458
rect 214760 477358 214788 597110
rect 216586 596728 216642 596737
rect 216586 596663 216642 596672
rect 214840 596488 214892 596494
rect 214840 596430 214892 596436
rect 214748 477352 214800 477358
rect 214748 477294 214800 477300
rect 214380 476342 214432 476348
rect 214654 476368 214710 476377
rect 214654 476303 214710 476312
rect 214760 476202 214788 477294
rect 214852 477290 214880 596430
rect 215116 596420 215168 596426
rect 215116 596362 215168 596368
rect 215024 596284 215076 596290
rect 215024 596226 215076 596232
rect 214932 563780 214984 563786
rect 214932 563722 214984 563728
rect 214840 477284 214892 477290
rect 214840 477226 214892 477232
rect 214852 476338 214880 477226
rect 214840 476332 214892 476338
rect 214840 476274 214892 476280
rect 214748 476196 214800 476202
rect 214748 476138 214800 476144
rect 214840 474428 214892 474434
rect 214840 474370 214892 474376
rect 214564 451920 214616 451926
rect 214564 451862 214616 451868
rect 214472 445324 214524 445330
rect 214472 445266 214524 445272
rect 214288 445256 214340 445262
rect 214288 445198 214340 445204
rect 213826 355600 213882 355609
rect 213826 355535 213882 355544
rect 213460 350532 213512 350538
rect 213460 350474 213512 350480
rect 213184 342236 213236 342242
rect 213184 342178 213236 342184
rect 213196 340950 213224 342178
rect 213184 340944 213236 340950
rect 213184 340886 213236 340892
rect 214196 327888 214248 327894
rect 214196 327830 214248 327836
rect 213090 293176 213146 293185
rect 213090 293111 213146 293120
rect 213104 279970 213132 293111
rect 213276 282872 213328 282878
rect 213276 282814 213328 282820
rect 213288 279970 213316 282814
rect 213642 282704 213698 282713
rect 213642 282639 213698 282648
rect 213656 279970 213684 282639
rect 214208 279970 214236 327830
rect 214300 285297 214328 445198
rect 214286 285288 214342 285297
rect 214286 285223 214342 285232
rect 214484 285161 214512 445266
rect 214470 285152 214526 285161
rect 214470 285087 214526 285096
rect 214576 279970 214604 451862
rect 214748 445188 214800 445194
rect 214748 445130 214800 445136
rect 214656 445120 214708 445126
rect 214656 445062 214708 445068
rect 214668 282334 214696 445062
rect 214760 285433 214788 445130
rect 214852 359242 214880 474370
rect 214840 359236 214892 359242
rect 214840 359178 214892 359184
rect 214746 285424 214802 285433
rect 214746 285359 214802 285368
rect 214656 282328 214708 282334
rect 214656 282270 214708 282276
rect 214944 279970 214972 563722
rect 215036 477086 215064 596226
rect 215128 477358 215156 596362
rect 216312 594788 216364 594794
rect 216312 594730 216364 594736
rect 215208 594176 215260 594182
rect 215208 594118 215260 594124
rect 215116 477352 215168 477358
rect 215116 477294 215168 477300
rect 215024 477080 215076 477086
rect 215024 477022 215076 477028
rect 215036 470594 215064 477022
rect 215128 476270 215156 477294
rect 215116 476264 215168 476270
rect 215116 476206 215168 476212
rect 215036 470566 215156 470594
rect 215024 445392 215076 445398
rect 215024 445334 215076 445340
rect 215036 285025 215064 445334
rect 215128 355706 215156 470566
rect 215220 359786 215248 594118
rect 216324 480254 216352 594730
rect 216496 593972 216548 593978
rect 216496 593914 216548 593920
rect 216324 480226 216444 480254
rect 216416 477154 216444 480226
rect 216508 477494 216536 593914
rect 216496 477488 216548 477494
rect 216496 477430 216548 477436
rect 216404 477148 216456 477154
rect 216404 477090 216456 477096
rect 216416 476882 216444 477090
rect 216404 476876 216456 476882
rect 216404 476818 216456 476824
rect 216416 476354 216444 476818
rect 216508 476474 216536 477430
rect 216496 476468 216548 476474
rect 216496 476410 216548 476416
rect 216416 476326 216536 476354
rect 216404 476196 216456 476202
rect 216404 476138 216456 476144
rect 215852 474700 215904 474706
rect 215852 474642 215904 474648
rect 215760 474224 215812 474230
rect 215760 474166 215812 474172
rect 215208 359780 215260 359786
rect 215208 359722 215260 359728
rect 215772 359582 215800 474166
rect 215760 359576 215812 359582
rect 215760 359518 215812 359524
rect 215864 358426 215892 474642
rect 215944 474564 215996 474570
rect 215944 474506 215996 474512
rect 215852 358420 215904 358426
rect 215852 358362 215904 358368
rect 215956 358358 215984 474506
rect 216126 474056 216182 474065
rect 216126 473991 216182 474000
rect 216036 473952 216088 473958
rect 216036 473894 216088 473900
rect 216048 358494 216076 473894
rect 216036 358488 216088 358494
rect 216036 358430 216088 358436
rect 215944 358352 215996 358358
rect 215944 358294 215996 358300
rect 216140 358086 216168 473991
rect 216220 473884 216272 473890
rect 216220 473826 216272 473832
rect 216232 358154 216260 473826
rect 216312 473816 216364 473822
rect 216312 473758 216364 473764
rect 216220 358148 216272 358154
rect 216220 358090 216272 358096
rect 216128 358080 216180 358086
rect 216128 358022 216180 358028
rect 216324 358018 216352 473758
rect 216312 358012 216364 358018
rect 216312 357954 216364 357960
rect 216416 355774 216444 476138
rect 216404 355768 216456 355774
rect 216404 355710 216456 355716
rect 215116 355700 215168 355706
rect 215116 355642 215168 355648
rect 216508 355502 216536 476326
rect 216600 358601 216628 596663
rect 217152 585818 217180 635831
rect 217140 585812 217192 585818
rect 217140 585754 217192 585760
rect 216770 516216 216826 516225
rect 216770 516151 216826 516160
rect 216680 479936 216732 479942
rect 216680 479878 216732 479884
rect 216692 479398 216720 479878
rect 216680 479392 216732 479398
rect 216680 479334 216732 479340
rect 216692 370025 216720 479334
rect 216784 454714 216812 516151
rect 217152 515953 217180 585754
rect 217244 563718 217272 636783
rect 217874 633720 217930 633729
rect 217874 633655 217930 633664
rect 217690 632768 217746 632777
rect 217690 632703 217746 632712
rect 217598 631000 217654 631009
rect 217598 630935 217654 630944
rect 217506 629912 217562 629921
rect 217506 629847 217562 629856
rect 217414 628144 217470 628153
rect 217414 628079 217470 628088
rect 217324 594652 217376 594658
rect 217324 594594 217376 594600
rect 217232 563712 217284 563718
rect 217232 563654 217284 563660
rect 217244 516905 217272 563654
rect 217230 516896 217286 516905
rect 217230 516831 217286 516840
rect 217244 516225 217272 516831
rect 217230 516216 217286 516225
rect 217230 516151 217286 516160
rect 216954 515944 217010 515953
rect 216954 515879 217010 515888
rect 217138 515944 217194 515953
rect 217138 515879 217194 515888
rect 216864 480004 216916 480010
rect 216864 479946 216916 479952
rect 216876 479534 216904 479946
rect 216864 479528 216916 479534
rect 216864 479470 216916 479476
rect 216772 454708 216824 454714
rect 216772 454650 216824 454656
rect 216876 390561 216904 479470
rect 216968 450838 216996 515879
rect 217046 513768 217102 513777
rect 217046 513703 217102 513712
rect 217060 480049 217088 513703
rect 217138 512816 217194 512825
rect 217138 512751 217194 512760
rect 217046 480040 217102 480049
rect 217046 479975 217102 479984
rect 217060 478961 217088 479975
rect 217152 479874 217180 512751
rect 217140 479868 217192 479874
rect 217140 479810 217192 479816
rect 217046 478952 217102 478961
rect 217046 478887 217102 478896
rect 217048 477488 217100 477494
rect 217048 477430 217100 477436
rect 217060 477222 217088 477430
rect 217048 477216 217100 477222
rect 217048 477158 217100 477164
rect 217048 476468 217100 476474
rect 217048 476410 217100 476416
rect 216956 450832 217008 450838
rect 216956 450774 217008 450780
rect 216954 391912 217010 391921
rect 216954 391847 217010 391856
rect 216968 391105 216996 391847
rect 216954 391096 217010 391105
rect 216954 391031 217010 391040
rect 216862 390552 216918 390561
rect 216862 390487 216918 390496
rect 216678 370016 216734 370025
rect 216678 369951 216734 369960
rect 216862 369880 216918 369889
rect 216862 369815 216918 369824
rect 216876 368393 216904 369815
rect 216862 368384 216918 368393
rect 216862 368319 216918 368328
rect 216968 358698 216996 391031
rect 216956 358692 217008 358698
rect 216956 358634 217008 358640
rect 216586 358592 216642 358601
rect 216586 358527 216642 358536
rect 216496 355496 216548 355502
rect 216496 355438 216548 355444
rect 215760 352572 215812 352578
rect 215760 352514 215812 352520
rect 215772 351830 215800 352514
rect 215760 351824 215812 351830
rect 215760 351766 215812 351772
rect 216404 351824 216456 351830
rect 216404 351766 216456 351772
rect 215300 330608 215352 330614
rect 215300 330550 215352 330556
rect 215022 285016 215078 285025
rect 215022 284951 215078 284960
rect 215312 279970 215340 330550
rect 215850 282840 215906 282849
rect 215850 282775 215906 282784
rect 216218 282840 216274 282849
rect 216218 282775 216274 282784
rect 215864 279970 215892 282775
rect 216232 279970 216260 282775
rect 211816 279942 212060 279970
rect 212368 279942 212428 279970
rect 212736 279942 212796 279970
rect 213104 279942 213164 279970
rect 213288 279942 213532 279970
rect 213656 279942 213900 279970
rect 214208 279942 214268 279970
rect 214576 279942 214636 279970
rect 214944 279942 215004 279970
rect 215312 279942 215372 279970
rect 215740 279942 215892 279970
rect 216108 279942 216260 279970
rect 216416 279970 216444 351766
rect 217060 349110 217088 476410
rect 217152 392873 217180 479810
rect 217232 478916 217284 478922
rect 217232 478858 217284 478864
rect 217138 392864 217194 392873
rect 217138 392799 217194 392808
rect 217244 391921 217272 478858
rect 217336 477494 217364 594594
rect 217428 508201 217456 628079
rect 217520 509969 217548 629847
rect 217612 511057 217640 630935
rect 217704 512825 217732 632703
rect 217782 610056 217838 610065
rect 217782 609991 217838 610000
rect 217690 512816 217746 512825
rect 217690 512751 217746 512760
rect 217598 511048 217654 511057
rect 217598 510983 217654 510992
rect 217506 509960 217562 509969
rect 217506 509895 217562 509904
rect 217414 508192 217470 508201
rect 217414 508127 217470 508136
rect 217428 479806 217456 508127
rect 217416 479800 217468 479806
rect 217416 479742 217468 479748
rect 217324 477488 217376 477494
rect 217324 477430 217376 477436
rect 217428 470594 217456 479742
rect 217520 479534 217548 509895
rect 217612 480078 217640 510983
rect 217796 489977 217824 609991
rect 217888 513777 217916 633655
rect 258078 599584 258134 599593
rect 258078 599519 258134 599528
rect 277306 599584 277362 599593
rect 277306 599519 277362 599528
rect 235998 597544 236054 597553
rect 235998 597479 236054 597488
rect 236182 597544 236238 597553
rect 236182 597479 236238 597488
rect 237378 597544 237434 597553
rect 237378 597479 237434 597488
rect 243082 597544 243138 597553
rect 243082 597479 243138 597488
rect 244278 597544 244334 597553
rect 244278 597479 244334 597488
rect 245474 597544 245530 597553
rect 245474 597479 245530 597488
rect 246486 597544 246542 597553
rect 246486 597479 246542 597488
rect 247038 597544 247094 597553
rect 247038 597479 247094 597488
rect 248418 597544 248474 597553
rect 248418 597479 248474 597488
rect 249798 597544 249854 597553
rect 249798 597479 249854 597488
rect 252098 597544 252154 597553
rect 252098 597479 252154 597488
rect 253478 597544 253534 597553
rect 253478 597479 253534 597488
rect 254582 597544 254638 597553
rect 254582 597479 254638 597488
rect 255410 597544 255466 597553
rect 255410 597479 255466 597488
rect 256698 597544 256754 597553
rect 256698 597479 256754 597488
rect 219990 597136 220046 597145
rect 219990 597071 220046 597080
rect 219716 597032 219768 597038
rect 219716 596974 219768 596980
rect 218888 596964 218940 596970
rect 218888 596906 218940 596912
rect 217968 596692 218020 596698
rect 217968 596634 218020 596640
rect 217874 513768 217930 513777
rect 217874 513703 217930 513712
rect 217782 489968 217838 489977
rect 217782 489903 217838 489912
rect 217600 480072 217652 480078
rect 217600 480014 217652 480020
rect 217508 479528 217560 479534
rect 217508 479470 217560 479476
rect 217612 478922 217640 480014
rect 217796 479398 217824 489903
rect 217784 479392 217836 479398
rect 217784 479334 217836 479340
rect 217600 478916 217652 478922
rect 217600 478858 217652 478864
rect 217980 477193 218008 596634
rect 218796 596556 218848 596562
rect 218796 596498 218848 596504
rect 218704 594720 218756 594726
rect 218704 594662 218756 594668
rect 218426 488064 218482 488073
rect 218426 487999 218482 488008
rect 218336 478984 218388 478990
rect 218336 478926 218388 478932
rect 217506 477184 217562 477193
rect 217506 477119 217562 477128
rect 217966 477184 218022 477193
rect 217966 477119 218022 477128
rect 217520 476649 217548 477119
rect 217968 477012 218020 477018
rect 217968 476954 218020 476960
rect 217506 476640 217562 476649
rect 217506 476575 217562 476584
rect 217784 476264 217836 476270
rect 217784 476206 217836 476212
rect 217428 470566 217548 470594
rect 217324 450832 217376 450838
rect 217324 450774 217376 450780
rect 217336 450566 217364 450774
rect 217324 450560 217376 450566
rect 217324 450502 217376 450508
rect 217336 396001 217364 450502
rect 217322 395992 217378 396001
rect 217322 395927 217378 395936
rect 217324 392080 217376 392086
rect 217324 392022 217376 392028
rect 217230 391912 217286 391921
rect 217230 391847 217286 391856
rect 217230 388240 217286 388249
rect 217230 388175 217286 388184
rect 217244 358766 217272 388175
rect 217336 359446 217364 392022
rect 217520 389174 217548 470566
rect 217692 454708 217744 454714
rect 217692 454650 217744 454656
rect 217704 396953 217732 454650
rect 217690 396944 217746 396953
rect 217690 396879 217746 396888
rect 217600 393372 217652 393378
rect 217600 393314 217652 393320
rect 217428 389146 217548 389174
rect 217428 388249 217456 389146
rect 217414 388240 217470 388249
rect 217414 388175 217470 388184
rect 217414 368112 217470 368121
rect 217414 368047 217470 368056
rect 217324 359440 217376 359446
rect 217324 359382 217376 359388
rect 217232 358760 217284 358766
rect 217232 358702 217284 358708
rect 217244 354674 217272 358702
rect 217324 358692 217376 358698
rect 217324 358634 217376 358640
rect 217152 354646 217272 354674
rect 217048 349104 217100 349110
rect 217048 349046 217100 349052
rect 216772 340876 216824 340882
rect 216772 340818 216824 340824
rect 216784 279970 216812 340818
rect 217152 279970 217180 354646
rect 217336 289270 217364 358634
rect 217428 355230 217456 368047
rect 217612 355570 217640 393314
rect 217600 355564 217652 355570
rect 217600 355506 217652 355512
rect 217416 355224 217468 355230
rect 217416 355166 217468 355172
rect 217508 291916 217560 291922
rect 217508 291858 217560 291864
rect 217324 289264 217376 289270
rect 217324 289206 217376 289212
rect 217520 279970 217548 291858
rect 217704 289202 217732 396879
rect 217796 355366 217824 476206
rect 217980 476134 218008 476954
rect 218060 476808 218112 476814
rect 218060 476750 218112 476756
rect 217968 476128 218020 476134
rect 217968 476070 218020 476076
rect 217874 390552 217930 390561
rect 217874 390487 217930 390496
rect 217888 390017 217916 390487
rect 217874 390008 217930 390017
rect 217874 389943 217930 389952
rect 217888 358630 217916 389943
rect 217876 358624 217928 358630
rect 217876 358566 217928 358572
rect 217784 355360 217836 355366
rect 217784 355302 217836 355308
rect 217692 289196 217744 289202
rect 217692 289138 217744 289144
rect 217888 288454 217916 358566
rect 217980 340882 218008 476070
rect 218072 393378 218100 476750
rect 218150 474736 218206 474745
rect 218150 474671 218206 474680
rect 218164 393961 218192 474671
rect 218150 393952 218206 393961
rect 218150 393887 218206 393896
rect 218060 393372 218112 393378
rect 218060 393314 218112 393320
rect 218348 358562 218376 478926
rect 218336 358556 218388 358562
rect 218336 358498 218388 358504
rect 218440 354006 218468 487999
rect 218716 476882 218744 594662
rect 218808 477018 218836 596498
rect 218900 477329 218928 596906
rect 219072 596896 219124 596902
rect 219072 596838 219124 596844
rect 218980 596760 219032 596766
rect 218980 596702 219032 596708
rect 218886 477320 218942 477329
rect 218886 477255 218942 477264
rect 218992 477057 219020 596702
rect 218978 477048 219034 477057
rect 218796 477012 218848 477018
rect 218978 476983 219034 476992
rect 218796 476954 218848 476960
rect 219084 476921 219112 596838
rect 219256 596828 219308 596834
rect 219256 596770 219308 596776
rect 219164 596624 219216 596630
rect 219164 596566 219216 596572
rect 219070 476912 219126 476921
rect 218704 476876 218756 476882
rect 219070 476847 219126 476856
rect 218704 476818 218756 476824
rect 219176 476746 219204 596566
rect 219268 477465 219296 596770
rect 219348 593904 219400 593910
rect 219348 593846 219400 593852
rect 219254 477456 219310 477465
rect 219254 477391 219310 477400
rect 219360 477222 219388 593846
rect 219728 478922 219756 596974
rect 219808 596352 219860 596358
rect 219808 596294 219860 596300
rect 219716 478916 219768 478922
rect 219716 478858 219768 478864
rect 219348 477216 219400 477222
rect 219348 477158 219400 477164
rect 219256 476876 219308 476882
rect 219256 476818 219308 476824
rect 219164 476740 219216 476746
rect 219164 476682 219216 476688
rect 219072 474632 219124 474638
rect 219072 474574 219124 474580
rect 218886 474192 218942 474201
rect 218704 474156 218756 474162
rect 218886 474127 218942 474136
rect 218704 474098 218756 474104
rect 218610 393816 218666 393825
rect 218610 393751 218666 393760
rect 218518 392864 218574 392873
rect 218518 392799 218574 392808
rect 218532 392018 218560 392799
rect 218520 392012 218572 392018
rect 218520 391954 218572 391960
rect 218518 368384 218574 368393
rect 218518 368319 218574 368328
rect 218532 359990 218560 368319
rect 218624 360058 218652 393751
rect 218716 392086 218744 474098
rect 218794 395992 218850 396001
rect 218794 395927 218850 395936
rect 218704 392080 218756 392086
rect 218704 392022 218756 392028
rect 218704 391944 218756 391950
rect 218704 391886 218756 391892
rect 218612 360052 218664 360058
rect 218612 359994 218664 360000
rect 218520 359984 218572 359990
rect 218520 359926 218572 359932
rect 218716 357950 218744 391886
rect 218704 357944 218756 357950
rect 218704 357886 218756 357892
rect 218808 355298 218836 395927
rect 218900 357882 218928 474127
rect 218980 446412 219032 446418
rect 218980 446354 219032 446360
rect 218888 357876 218940 357882
rect 218888 357818 218940 357824
rect 218796 355292 218848 355298
rect 218796 355234 218848 355240
rect 218428 354000 218480 354006
rect 218428 353942 218480 353948
rect 217968 340876 218020 340882
rect 217968 340818 218020 340824
rect 218612 293820 218664 293826
rect 218612 293762 218664 293768
rect 217876 288448 217928 288454
rect 217876 288390 217928 288396
rect 217690 282840 217746 282849
rect 217690 282775 217746 282784
rect 218426 282840 218482 282849
rect 218426 282775 218482 282784
rect 217704 279970 217732 282775
rect 218440 279970 218468 282775
rect 216416 279942 216476 279970
rect 216784 279942 216844 279970
rect 217152 279942 217212 279970
rect 217520 279942 217580 279970
rect 217704 279942 217948 279970
rect 218316 279942 218468 279970
rect 218624 279970 218652 293762
rect 218992 279970 219020 446354
rect 219084 358290 219112 474574
rect 219072 358284 219124 358290
rect 219072 358226 219124 358232
rect 219268 355434 219296 476818
rect 219360 476814 219388 477158
rect 219348 476808 219400 476814
rect 219348 476750 219400 476756
rect 219820 476542 219848 596294
rect 219900 594380 219952 594386
rect 219900 594322 219952 594328
rect 219808 476536 219860 476542
rect 219808 476478 219860 476484
rect 219716 474496 219768 474502
rect 219716 474438 219768 474444
rect 219624 474360 219676 474366
rect 219624 474302 219676 474308
rect 219636 359378 219664 474302
rect 219624 359372 219676 359378
rect 219624 359314 219676 359320
rect 219346 358456 219402 358465
rect 219346 358391 219402 358400
rect 219256 355428 219308 355434
rect 219256 355370 219308 355376
rect 219360 279970 219388 358391
rect 219728 358222 219756 474438
rect 219716 358216 219768 358222
rect 219716 358158 219768 358164
rect 219820 353258 219848 476478
rect 219912 474745 219940 594322
rect 219898 474736 219954 474745
rect 219898 474671 219954 474680
rect 219900 443692 219952 443698
rect 219900 443634 219952 443640
rect 219808 353252 219860 353258
rect 219808 353194 219860 353200
rect 219716 297424 219768 297430
rect 219716 297366 219768 297372
rect 219728 279970 219756 297366
rect 219912 282878 219940 443634
rect 220004 358057 220032 597071
rect 236012 597038 236040 597479
rect 236000 597032 236052 597038
rect 236000 596974 236052 596980
rect 236196 596970 236224 597479
rect 236184 596964 236236 596970
rect 236184 596906 236236 596912
rect 237392 596902 237420 597479
rect 243096 597106 243124 597479
rect 243084 597100 243136 597106
rect 243084 597042 243136 597048
rect 237380 596896 237432 596902
rect 237380 596838 237432 596844
rect 238758 596864 238814 596873
rect 238758 596799 238760 596808
rect 238812 596799 238814 596808
rect 240138 596864 240194 596873
rect 240138 596799 240194 596808
rect 241518 596864 241574 596873
rect 241518 596799 241574 596808
rect 238760 596770 238812 596776
rect 240152 596766 240180 596799
rect 240140 596760 240192 596766
rect 240140 596702 240192 596708
rect 241532 596698 241560 596799
rect 241520 596692 241572 596698
rect 241520 596634 241572 596640
rect 243096 596630 243124 597042
rect 244292 597038 244320 597479
rect 244280 597032 244332 597038
rect 244280 596974 244332 596980
rect 243084 596624 243136 596630
rect 243084 596566 243136 596572
rect 244292 596562 244320 596974
rect 245488 596970 245516 597479
rect 244372 596964 244424 596970
rect 244372 596906 244424 596912
rect 245476 596964 245528 596970
rect 245476 596906 245528 596912
rect 244280 596556 244332 596562
rect 244280 596498 244332 596504
rect 244384 596494 244412 596906
rect 246500 596834 246528 597479
rect 245660 596828 245712 596834
rect 245660 596770 245712 596776
rect 246488 596828 246540 596834
rect 246488 596770 246540 596776
rect 244372 596488 244424 596494
rect 244372 596430 244424 596436
rect 245672 596426 245700 596770
rect 245660 596420 245712 596426
rect 245660 596362 245712 596368
rect 247052 566545 247080 597479
rect 247130 596864 247186 596873
rect 247130 596799 247186 596808
rect 247144 596494 247172 596799
rect 248432 596630 248460 597479
rect 248420 596624 248472 596630
rect 248420 596566 248472 596572
rect 247132 596488 247184 596494
rect 247132 596430 247184 596436
rect 247144 594046 247172 596430
rect 247132 594040 247184 594046
rect 247132 593982 247184 593988
rect 248432 593978 248460 596566
rect 248420 593972 248472 593978
rect 248420 593914 248472 593920
rect 247038 566536 247094 566545
rect 247038 566471 247094 566480
rect 249812 563786 249840 597479
rect 249890 596864 249946 596873
rect 249890 596799 249946 596808
rect 249904 596562 249932 596799
rect 252112 596766 252140 597479
rect 252190 596864 252246 596873
rect 252190 596799 252246 596808
rect 252100 596760 252152 596766
rect 252100 596702 252152 596708
rect 249892 596556 249944 596562
rect 249892 596498 249944 596504
rect 249904 594794 249932 596498
rect 249892 594788 249944 594794
rect 249892 594730 249944 594736
rect 252112 594658 252140 596702
rect 252204 596698 252232 596799
rect 252192 596692 252244 596698
rect 252192 596634 252244 596640
rect 252100 594652 252152 594658
rect 252100 594594 252152 594600
rect 252204 593910 252232 596634
rect 253492 596426 253520 597479
rect 254596 596902 254624 597479
rect 253940 596896 253992 596902
rect 253940 596838 253992 596844
rect 254584 596896 254636 596902
rect 254584 596838 254636 596844
rect 253480 596420 253532 596426
rect 253480 596362 253532 596368
rect 253492 594726 253520 596362
rect 253952 596358 253980 596838
rect 253940 596352 253992 596358
rect 253940 596294 253992 596300
rect 255424 596222 255452 597479
rect 256712 597242 256740 597479
rect 256700 597236 256752 597242
rect 256700 597178 256752 597184
rect 256712 596290 256740 597178
rect 258092 597174 258120 599519
rect 260838 597544 260894 597553
rect 260838 597479 260894 597488
rect 263598 597544 263654 597553
rect 263598 597479 263654 597488
rect 264978 597544 265034 597553
rect 264978 597479 265034 597488
rect 267738 597544 267794 597553
rect 267738 597479 267794 597488
rect 270498 597544 270554 597553
rect 270498 597479 270554 597488
rect 276018 597544 276074 597553
rect 276018 597479 276074 597488
rect 258080 597168 258132 597174
rect 258080 597110 258132 597116
rect 260852 597106 260880 597479
rect 262218 597408 262274 597417
rect 262218 597343 262274 597352
rect 260840 597100 260892 597106
rect 260840 597042 260892 597048
rect 262232 597038 262260 597343
rect 262220 597032 262272 597038
rect 262220 596974 262272 596980
rect 259550 596728 259606 596737
rect 259550 596663 259606 596672
rect 259458 596592 259514 596601
rect 259458 596527 259514 596536
rect 256700 596284 256752 596290
rect 256700 596226 256752 596232
rect 255412 596216 255464 596222
rect 255412 596158 255464 596164
rect 253480 594720 253532 594726
rect 253480 594662 253532 594668
rect 255424 594590 255452 596158
rect 255412 594584 255464 594590
rect 255412 594526 255464 594532
rect 259472 594522 259500 596527
rect 259460 594516 259512 594522
rect 259460 594458 259512 594464
rect 259564 594454 259592 596663
rect 263612 594561 263640 597479
rect 263690 597408 263746 597417
rect 263690 597343 263746 597352
rect 263704 596970 263732 597343
rect 263692 596964 263744 596970
rect 263692 596906 263744 596912
rect 263598 594552 263654 594561
rect 263598 594487 263654 594496
rect 259552 594448 259604 594454
rect 264992 594425 265020 597479
rect 266358 597408 266414 597417
rect 266358 597343 266414 597352
rect 265070 596864 265126 596873
rect 265070 596799 265072 596808
rect 265124 596799 265126 596808
rect 265072 596770 265124 596776
rect 266372 596630 266400 597343
rect 266360 596624 266412 596630
rect 266360 596566 266412 596572
rect 266360 596488 266412 596494
rect 266358 596456 266360 596465
rect 266412 596456 266414 596465
rect 266358 596391 266414 596400
rect 259552 594390 259604 594396
rect 264978 594416 265034 594425
rect 264978 594351 265034 594360
rect 267752 594289 267780 597479
rect 270406 597408 270462 597417
rect 270406 597343 270462 597352
rect 270420 597145 270448 597343
rect 270406 597136 270462 597145
rect 270406 597071 270462 597080
rect 267922 596728 267978 596737
rect 267922 596663 267978 596672
rect 269118 596728 269174 596737
rect 269118 596663 269120 596672
rect 267936 596562 267964 596663
rect 269172 596663 269174 596672
rect 269120 596634 269172 596640
rect 267924 596556 267976 596562
rect 267924 596498 267976 596504
rect 267738 594280 267794 594289
rect 267738 594215 267794 594224
rect 270512 594153 270540 597479
rect 274638 597272 274694 597281
rect 274638 597207 274640 597216
rect 274692 597207 274694 597216
rect 274640 597178 274692 597184
rect 276032 597174 276060 597479
rect 276020 597168 276072 597174
rect 270590 597136 270646 597145
rect 270590 597071 270646 597080
rect 273258 597136 273314 597145
rect 276020 597110 276072 597116
rect 273258 597071 273314 597080
rect 270604 596766 270632 597071
rect 273272 596902 273300 597071
rect 277320 597009 277348 599519
rect 280158 597544 280214 597553
rect 280158 597479 280214 597488
rect 282918 597544 282974 597553
rect 282918 597479 282974 597488
rect 285678 597544 285734 597553
rect 285678 597479 285734 597488
rect 289818 597544 289874 597553
rect 289818 597479 289874 597488
rect 292578 597544 292634 597553
rect 292578 597479 292634 597488
rect 277306 597000 277362 597009
rect 277306 596935 277362 596944
rect 273260 596896 273312 596902
rect 273260 596838 273312 596844
rect 270592 596760 270644 596766
rect 270592 596702 270644 596708
rect 271878 596456 271934 596465
rect 271878 596391 271880 596400
rect 271932 596391 271934 596400
rect 271880 596362 271932 596368
rect 273258 596320 273314 596329
rect 273258 596255 273314 596264
rect 273272 596222 273300 596255
rect 273260 596216 273312 596222
rect 273260 596158 273312 596164
rect 280172 594318 280200 597479
rect 280160 594312 280212 594318
rect 280160 594254 280212 594260
rect 270498 594144 270554 594153
rect 270498 594079 270554 594088
rect 282932 594017 282960 597479
rect 285692 594386 285720 597479
rect 287058 597136 287114 597145
rect 287058 597071 287114 597080
rect 285680 594380 285732 594386
rect 285680 594322 285732 594328
rect 287072 594250 287100 597071
rect 287060 594244 287112 594250
rect 287060 594186 287112 594192
rect 289832 594114 289860 597479
rect 292592 594182 292620 597479
rect 326986 597000 327042 597009
rect 326986 596935 327042 596944
rect 327000 596902 327028 596935
rect 326988 596896 327040 596902
rect 311806 596864 311862 596873
rect 311806 596799 311862 596808
rect 321466 596864 321522 596873
rect 321466 596799 321522 596808
rect 324226 596864 324282 596873
rect 326988 596838 327040 596844
rect 356794 596864 356850 596873
rect 324226 596799 324228 596808
rect 311820 596494 311848 596799
rect 321480 596766 321508 596799
rect 324280 596799 324282 596808
rect 356794 596799 356850 596808
rect 357900 596828 357952 596834
rect 324228 596770 324280 596776
rect 321468 596760 321520 596766
rect 314566 596728 314622 596737
rect 314566 596663 314622 596672
rect 318706 596728 318762 596737
rect 321468 596702 321520 596708
rect 318706 596663 318708 596672
rect 314580 596630 314608 596663
rect 318760 596663 318762 596672
rect 318708 596634 318760 596640
rect 314568 596624 314620 596630
rect 314568 596566 314620 596572
rect 315946 596592 316002 596601
rect 315946 596527 315948 596536
rect 316000 596527 316002 596536
rect 315948 596498 316000 596504
rect 311808 596488 311860 596494
rect 306102 596456 306158 596465
rect 306102 596391 306158 596400
rect 309046 596456 309102 596465
rect 311808 596430 311860 596436
rect 309046 596391 309048 596400
rect 306116 596358 306144 596391
rect 309100 596391 309102 596400
rect 356612 596420 356664 596426
rect 309048 596362 309100 596368
rect 356612 596362 356664 596368
rect 306104 596352 306156 596358
rect 296350 596320 296406 596329
rect 296350 596255 296406 596264
rect 303526 596320 303582 596329
rect 306104 596294 306156 596300
rect 303526 596255 303528 596264
rect 296364 596222 296392 596255
rect 303580 596255 303582 596264
rect 303528 596226 303580 596232
rect 296352 596216 296404 596222
rect 296352 596158 296404 596164
rect 292580 594176 292632 594182
rect 292580 594118 292632 594124
rect 289820 594108 289872 594114
rect 289820 594050 289872 594056
rect 282918 594008 282974 594017
rect 282918 593943 282974 593952
rect 252192 593904 252244 593910
rect 252192 593846 252244 593852
rect 351092 567180 351144 567186
rect 351092 567122 351144 567128
rect 351104 565865 351132 567122
rect 351090 565856 351146 565865
rect 351090 565791 351146 565800
rect 249800 563780 249852 563786
rect 249800 563722 249852 563728
rect 235998 479632 236054 479641
rect 235998 479567 236054 479576
rect 236012 478922 236040 479567
rect 236000 478916 236052 478922
rect 236000 478858 236052 478864
rect 252376 477488 252428 477494
rect 243174 477456 243230 477465
rect 243174 477391 243230 477400
rect 244278 477456 244334 477465
rect 244278 477391 244334 477400
rect 245474 477456 245530 477465
rect 245474 477391 245530 477400
rect 245934 477456 245990 477465
rect 245934 477391 245990 477400
rect 247130 477456 247186 477465
rect 247130 477391 247186 477400
rect 248602 477456 248658 477465
rect 248602 477391 248658 477400
rect 250074 477456 250130 477465
rect 250074 477391 250130 477400
rect 251270 477456 251326 477465
rect 251270 477391 251326 477400
rect 252374 477456 252376 477465
rect 252468 477488 252520 477494
rect 252428 477456 252430 477465
rect 269120 477488 269172 477494
rect 252468 477430 252520 477436
rect 253386 477456 253442 477465
rect 252374 477391 252430 477400
rect 220728 476808 220780 476814
rect 220728 476750 220780 476756
rect 220740 476542 220768 476750
rect 243188 476746 243216 477391
rect 244292 477018 244320 477391
rect 245488 477290 245516 477391
rect 245948 477358 245976 477391
rect 247144 477358 247172 477391
rect 245936 477352 245988 477358
rect 245936 477294 245988 477300
rect 247132 477352 247184 477358
rect 247132 477294 247184 477300
rect 245476 477284 245528 477290
rect 245476 477226 245528 477232
rect 244280 477012 244332 477018
rect 244280 476954 244332 476960
rect 243176 476740 243228 476746
rect 243176 476682 243228 476688
rect 244292 476542 244320 476954
rect 245948 476950 245976 477294
rect 245936 476944 245988 476950
rect 245936 476886 245988 476892
rect 220728 476536 220780 476542
rect 220728 476478 220780 476484
rect 244280 476536 244332 476542
rect 244280 476478 244332 476484
rect 247144 476270 247172 477294
rect 248616 476678 248644 477391
rect 250088 477154 250116 477391
rect 251284 477222 251312 477391
rect 251272 477216 251324 477222
rect 251272 477158 251324 477164
rect 250076 477148 250128 477154
rect 250076 477090 250128 477096
rect 251088 477148 251140 477154
rect 251088 477090 251140 477096
rect 248604 476672 248656 476678
rect 248604 476614 248656 476620
rect 251100 476610 251128 477090
rect 252388 477018 252416 477391
rect 252480 477222 252508 477430
rect 253386 477391 253442 477400
rect 254490 477456 254546 477465
rect 254490 477391 254546 477400
rect 255318 477456 255374 477465
rect 255318 477391 255320 477400
rect 252468 477216 252520 477222
rect 252468 477158 252520 477164
rect 252376 477012 252428 477018
rect 252376 476954 252428 476960
rect 253400 476882 253428 477391
rect 253388 476876 253440 476882
rect 253388 476818 253440 476824
rect 254504 476814 254532 477391
rect 255372 477391 255374 477400
rect 256974 477456 257030 477465
rect 256974 477391 257030 477400
rect 260838 477456 260894 477465
rect 260838 477391 260840 477400
rect 255320 477362 255372 477368
rect 255332 477154 255360 477362
rect 255320 477148 255372 477154
rect 255320 477090 255372 477096
rect 256988 477086 257016 477391
rect 260892 477391 260894 477400
rect 266358 477456 266414 477465
rect 266358 477391 266414 477400
rect 269118 477456 269120 477465
rect 269172 477456 269174 477465
rect 269118 477391 269174 477400
rect 278778 477456 278834 477465
rect 278778 477391 278780 477400
rect 260840 477362 260892 477368
rect 266372 477358 266400 477391
rect 278832 477391 278834 477400
rect 278780 477362 278832 477368
rect 266360 477352 266412 477358
rect 259366 477320 259422 477329
rect 259366 477255 259422 477264
rect 260838 477320 260894 477329
rect 260838 477255 260894 477264
rect 263598 477320 263654 477329
rect 266360 477294 266412 477300
rect 271878 477320 271934 477329
rect 263598 477255 263600 477264
rect 259380 477222 259408 477255
rect 259368 477216 259420 477222
rect 259368 477158 259420 477164
rect 256976 477080 257028 477086
rect 256976 477022 257028 477028
rect 255318 476912 255374 476921
rect 255318 476847 255374 476856
rect 254492 476808 254544 476814
rect 254492 476750 254544 476756
rect 251088 476604 251140 476610
rect 251088 476546 251140 476552
rect 247132 476264 247184 476270
rect 247038 476232 247094 476241
rect 247132 476206 247184 476212
rect 249798 476232 249854 476241
rect 247038 476167 247094 476176
rect 249798 476167 249854 476176
rect 252558 476232 252614 476241
rect 252558 476167 252614 476176
rect 247052 449274 247080 476167
rect 249812 451926 249840 476167
rect 249800 451920 249852 451926
rect 249800 451862 249852 451868
rect 247040 449268 247092 449274
rect 247040 449210 247092 449216
rect 252572 446418 252600 476167
rect 255332 474201 255360 476847
rect 258262 476232 258318 476241
rect 259380 476202 259408 477158
rect 260852 476746 260880 477255
rect 263652 477255 263654 477264
rect 263692 477284 263744 477290
rect 263600 477226 263652 477232
rect 271878 477255 271934 477264
rect 276018 477320 276074 477329
rect 276018 477255 276074 477264
rect 277674 477320 277730 477329
rect 277674 477255 277676 477264
rect 263692 477226 263744 477232
rect 262218 476912 262274 476921
rect 262218 476847 262274 476856
rect 260840 476740 260892 476746
rect 260840 476682 260892 476688
rect 262232 476542 262260 476847
rect 263704 476649 263732 477226
rect 264978 477048 265034 477057
rect 264978 476983 265034 476992
rect 270498 477048 270554 477057
rect 270498 476983 270500 476992
rect 264992 476950 265020 476983
rect 270552 476983 270554 476992
rect 270500 476954 270552 476960
rect 264980 476944 265032 476950
rect 264980 476886 265032 476892
rect 270498 476912 270554 476921
rect 271892 476882 271920 477255
rect 276032 477222 276060 477255
rect 277728 477255 277730 477264
rect 277676 477226 277728 477232
rect 276020 477216 276072 477222
rect 273258 477184 273314 477193
rect 273258 477119 273260 477128
rect 273312 477119 273314 477128
rect 274638 477184 274694 477193
rect 276020 477158 276072 477164
rect 311806 477184 311862 477193
rect 274638 477119 274694 477128
rect 311806 477119 311862 477128
rect 273260 477090 273312 477096
rect 274652 477086 274680 477119
rect 274640 477080 274692 477086
rect 274640 477022 274692 477028
rect 277582 477048 277638 477057
rect 277582 476983 277638 476992
rect 285678 477048 285734 477057
rect 285678 476983 285734 476992
rect 273258 476912 273314 476921
rect 270498 476847 270554 476856
rect 271880 476876 271932 476882
rect 266358 476776 266414 476785
rect 266358 476711 266414 476720
rect 266372 476678 266400 476711
rect 266360 476672 266412 476678
rect 263690 476640 263746 476649
rect 266360 476614 266412 476620
rect 268198 476640 268254 476649
rect 263690 476575 263746 476584
rect 268198 476575 268200 476584
rect 268252 476575 268254 476584
rect 268200 476546 268252 476552
rect 262220 476536 262272 476542
rect 262220 476478 262272 476484
rect 260838 476232 260894 476241
rect 258262 476167 258318 476176
rect 259368 476196 259420 476202
rect 255318 474192 255374 474201
rect 255318 474127 255374 474136
rect 258276 474065 258304 476167
rect 260838 476167 260894 476176
rect 263598 476232 263654 476241
rect 263598 476167 263654 476176
rect 264978 476232 265034 476241
rect 264978 476167 265034 476176
rect 268014 476232 268070 476241
rect 268014 476167 268070 476176
rect 259368 476138 259420 476144
rect 258262 474056 258318 474065
rect 258262 473991 258318 474000
rect 260852 473822 260880 476167
rect 263612 473890 263640 476167
rect 264992 473958 265020 476167
rect 268028 474706 268056 476167
rect 268016 474700 268068 474706
rect 268016 474642 268068 474648
rect 270512 474570 270540 476847
rect 273258 476847 273314 476856
rect 271880 476818 271932 476824
rect 273272 476814 273300 476847
rect 273260 476808 273312 476814
rect 273260 476750 273312 476756
rect 273258 476232 273314 476241
rect 273258 476167 273314 476176
rect 276018 476232 276074 476241
rect 276018 476167 276074 476176
rect 273272 474638 273300 476167
rect 273260 474632 273312 474638
rect 273260 474574 273312 474580
rect 270500 474564 270552 474570
rect 270500 474506 270552 474512
rect 276032 474502 276060 476167
rect 276020 474496 276072 474502
rect 276020 474438 276072 474444
rect 277596 474434 277624 476983
rect 280158 476232 280214 476241
rect 280158 476167 280214 476176
rect 282918 476232 282974 476241
rect 282918 476167 282974 476176
rect 277584 474428 277636 474434
rect 277584 474370 277636 474376
rect 280172 474298 280200 476167
rect 280160 474292 280212 474298
rect 280160 474234 280212 474240
rect 282932 474230 282960 476167
rect 285692 474366 285720 476983
rect 287702 476776 287758 476785
rect 287702 476711 287758 476720
rect 302146 476776 302202 476785
rect 302146 476711 302202 476720
rect 285680 474360 285732 474366
rect 285680 474302 285732 474308
rect 282920 474224 282972 474230
rect 282920 474166 282972 474172
rect 287716 474094 287744 476711
rect 289818 476504 289874 476513
rect 289818 476439 289874 476448
rect 287704 474088 287756 474094
rect 287704 474030 287756 474036
rect 289832 474026 289860 476439
rect 299386 476368 299442 476377
rect 299386 476303 299442 476312
rect 292578 476232 292634 476241
rect 292578 476167 292634 476176
rect 296258 476232 296314 476241
rect 299400 476202 299428 476303
rect 302160 476270 302188 476711
rect 309046 476640 309102 476649
rect 309046 476575 309102 476584
rect 306102 476504 306158 476513
rect 309060 476474 309088 476575
rect 311820 476542 311848 477119
rect 324226 477048 324282 477057
rect 324226 476983 324282 476992
rect 326986 477048 327042 477057
rect 326986 476983 327042 476992
rect 321466 476912 321522 476921
rect 324240 476882 324268 476983
rect 327000 476950 327028 476983
rect 326988 476944 327040 476950
rect 326988 476886 327040 476892
rect 321466 476847 321522 476856
rect 324228 476876 324280 476882
rect 321480 476814 321508 476847
rect 324228 476818 324280 476824
rect 321468 476808 321520 476814
rect 315946 476776 316002 476785
rect 315946 476711 316002 476720
rect 318706 476776 318762 476785
rect 321468 476750 321520 476756
rect 318706 476711 318708 476720
rect 315960 476678 315988 476711
rect 318760 476711 318762 476720
rect 318708 476682 318760 476688
rect 315948 476672 316000 476678
rect 314566 476640 314622 476649
rect 315948 476614 316000 476620
rect 314566 476575 314568 476584
rect 314620 476575 314622 476584
rect 314568 476546 314620 476552
rect 311808 476536 311860 476542
rect 311808 476478 311860 476484
rect 306102 476439 306158 476448
rect 309048 476468 309100 476474
rect 306116 476406 306144 476439
rect 309048 476410 309100 476416
rect 306104 476400 306156 476406
rect 303526 476368 303582 476377
rect 306104 476342 306156 476348
rect 303526 476303 303528 476312
rect 303580 476303 303582 476312
rect 303528 476274 303580 476280
rect 302148 476264 302200 476270
rect 302148 476206 302200 476212
rect 296258 476167 296314 476176
rect 299388 476196 299440 476202
rect 292592 474162 292620 476167
rect 296272 476134 296300 476167
rect 299388 476138 299440 476144
rect 296260 476128 296312 476134
rect 296260 476070 296312 476076
rect 292580 474156 292632 474162
rect 292580 474098 292632 474104
rect 289820 474020 289872 474026
rect 289820 473962 289872 473968
rect 264980 473952 265032 473958
rect 264980 473894 265032 473900
rect 263600 473884 263652 473890
rect 263600 473826 263652 473832
rect 260840 473816 260892 473822
rect 260840 473758 260892 473764
rect 351092 447092 351144 447098
rect 351092 447034 351144 447040
rect 252560 446412 252612 446418
rect 252560 446354 252612 446360
rect 351104 445777 351132 447034
rect 351090 445768 351146 445777
rect 351090 445703 351146 445712
rect 224224 360052 224276 360058
rect 224224 359994 224276 360000
rect 234068 360052 234120 360058
rect 234068 359994 234120 360000
rect 221922 359952 221978 359961
rect 221922 359887 221978 359896
rect 219990 358048 220046 358057
rect 219990 357983 220046 357992
rect 220082 311128 220138 311137
rect 220082 311063 220138 311072
rect 219900 282872 219952 282878
rect 219900 282814 219952 282820
rect 220096 279970 220124 311063
rect 221556 288448 221608 288454
rect 221556 288390 221608 288396
rect 220820 287972 220872 287978
rect 220820 287914 220872 287920
rect 220266 282840 220322 282849
rect 220266 282775 220322 282784
rect 220280 279970 220308 282775
rect 220832 279970 220860 287914
rect 221464 286544 221516 286550
rect 221464 286486 221516 286492
rect 221476 279970 221504 286486
rect 218624 279942 218684 279970
rect 218992 279942 219052 279970
rect 219360 279942 219420 279970
rect 219728 279942 219788 279970
rect 220096 279942 220156 279970
rect 220280 279942 220524 279970
rect 220832 279942 220892 279970
rect 221260 279942 221504 279970
rect 221568 279970 221596 288390
rect 221936 279970 221964 359887
rect 223762 358728 223818 358737
rect 223762 358663 223818 358672
rect 223396 357876 223448 357882
rect 223396 357818 223448 357824
rect 223028 330676 223080 330682
rect 223028 330618 223080 330624
rect 222476 285252 222528 285258
rect 222476 285194 222528 285200
rect 222200 282872 222252 282878
rect 222200 282814 222252 282820
rect 222212 279970 222240 282814
rect 222488 279970 222516 285194
rect 223040 279970 223068 330618
rect 223408 279970 223436 357818
rect 223776 279970 223804 358663
rect 224236 358465 224264 359994
rect 228178 358592 228234 358601
rect 228178 358527 228234 358536
rect 224222 358456 224278 358465
rect 224222 358391 224278 358400
rect 227812 358080 227864 358086
rect 227812 358022 227864 358028
rect 225234 356688 225290 356697
rect 225234 356623 225290 356632
rect 225248 355162 225276 356623
rect 225236 355156 225288 355162
rect 225236 355098 225288 355104
rect 224868 337476 224920 337482
rect 224868 337418 224920 337424
rect 224132 331900 224184 331906
rect 224132 331842 224184 331848
rect 224144 279970 224172 331842
rect 224500 312588 224552 312594
rect 224500 312530 224552 312536
rect 224512 279970 224540 312530
rect 224880 279970 224908 337418
rect 225248 279970 225276 355098
rect 226340 354000 226392 354006
rect 226340 353942 226392 353948
rect 225328 351348 225380 351354
rect 225328 351290 225380 351296
rect 225340 350538 225368 351290
rect 225328 350532 225380 350538
rect 225328 350474 225380 350480
rect 225604 350532 225656 350538
rect 225604 350474 225656 350480
rect 225616 279970 225644 350474
rect 225972 289264 226024 289270
rect 225972 289206 226024 289212
rect 225984 279970 226012 289206
rect 226352 279970 226380 353942
rect 227444 340264 227496 340270
rect 227444 340206 227496 340212
rect 227074 291000 227130 291009
rect 227074 290935 227130 290944
rect 226524 282396 226576 282402
rect 226524 282338 226576 282344
rect 226536 279970 226564 282338
rect 227088 279970 227116 290935
rect 227456 279970 227484 340206
rect 227824 279970 227852 358022
rect 228192 279970 228220 358527
rect 234080 358465 234108 359994
rect 270500 359916 270552 359922
rect 270500 359858 270552 359864
rect 311716 359916 311768 359922
rect 311716 359858 311768 359864
rect 263874 359680 263930 359689
rect 263874 359615 263930 359624
rect 270132 359644 270184 359650
rect 263508 359576 263560 359582
rect 253202 359544 253258 359553
rect 263508 359518 263560 359524
rect 253202 359479 253258 359488
rect 259736 359508 259788 359514
rect 253216 359281 253244 359479
rect 259736 359450 259788 359456
rect 261300 359508 261352 359514
rect 261300 359450 261352 359456
rect 257252 359304 257304 359310
rect 253202 359272 253258 359281
rect 257252 359246 257304 359252
rect 253202 359207 253258 359216
rect 256884 359236 256936 359242
rect 256884 359178 256936 359184
rect 235998 358592 236054 358601
rect 235998 358527 236000 358536
rect 236052 358527 236054 358536
rect 236000 358498 236052 358504
rect 234066 358456 234122 358465
rect 234066 358391 234122 358400
rect 232226 358320 232282 358329
rect 232226 358255 232282 358264
rect 231860 358012 231912 358018
rect 231860 357954 231912 357960
rect 230020 357944 230072 357950
rect 230020 357886 230072 357892
rect 228548 342916 228600 342922
rect 228548 342858 228600 342864
rect 228560 279970 228588 342858
rect 229282 298752 229338 298761
rect 229282 298687 229338 298696
rect 228916 297560 228968 297566
rect 228916 297502 228968 297508
rect 228928 279970 228956 297502
rect 229296 279970 229324 298687
rect 229928 285252 229980 285258
rect 229928 285194 229980 285200
rect 229940 279970 229968 285194
rect 221568 279942 221628 279970
rect 221936 279942 221996 279970
rect 222212 279942 222364 279970
rect 222488 279942 222732 279970
rect 223040 279942 223100 279970
rect 223408 279942 223468 279970
rect 223776 279942 223836 279970
rect 224144 279942 224204 279970
rect 224512 279942 224572 279970
rect 224880 279942 224940 279970
rect 225248 279942 225308 279970
rect 225616 279942 225676 279970
rect 225984 279942 226044 279970
rect 226352 279942 226412 279970
rect 226536 279942 226780 279970
rect 227088 279942 227148 279970
rect 227456 279942 227516 279970
rect 227824 279942 227884 279970
rect 228192 279942 228252 279970
rect 228560 279942 228620 279970
rect 228928 279942 228988 279970
rect 229296 279942 229356 279970
rect 229724 279942 229968 279970
rect 230032 279970 230060 357886
rect 230388 355224 230440 355230
rect 230388 355166 230440 355172
rect 230400 279970 230428 355166
rect 231492 354000 231544 354006
rect 231492 353942 231544 353948
rect 231124 293956 231176 293962
rect 231124 293898 231176 293904
rect 230572 285184 230624 285190
rect 230572 285126 230624 285132
rect 230584 279970 230612 285126
rect 231136 279970 231164 293898
rect 231504 279970 231532 353942
rect 231872 279970 231900 357954
rect 232240 279970 232268 358255
rect 233700 356176 233752 356182
rect 233700 356118 233752 356124
rect 233712 349110 233740 356118
rect 233700 349104 233752 349110
rect 233700 349046 233752 349052
rect 232596 327820 232648 327826
rect 232596 327762 232648 327768
rect 232608 279970 232636 327762
rect 232964 297628 233016 297634
rect 232964 297570 233016 297576
rect 232976 279970 233004 297570
rect 233330 297392 233386 297401
rect 233330 297327 233386 297336
rect 233344 279970 233372 297327
rect 233712 279970 233740 349046
rect 234080 279970 234108 358391
rect 236012 358154 236040 358498
rect 239956 358488 240008 358494
rect 239956 358430 240008 358436
rect 235908 358148 235960 358154
rect 235908 358090 235960 358096
rect 236000 358148 236052 358154
rect 236000 358090 236052 358096
rect 234434 325000 234490 325009
rect 234434 324935 234490 324944
rect 234448 279970 234476 324935
rect 235540 304360 235592 304366
rect 235540 304302 235592 304308
rect 235172 293888 235224 293894
rect 235172 293830 235224 293836
rect 234804 287904 234856 287910
rect 234804 287846 234856 287852
rect 234816 279970 234844 287846
rect 235184 279970 235212 293830
rect 235552 279970 235580 304302
rect 235920 279970 235948 358090
rect 236012 354674 236040 358090
rect 238022 357232 238078 357241
rect 238022 357167 238078 357176
rect 237010 356280 237066 356289
rect 237010 356215 237066 356224
rect 236274 355872 236330 355881
rect 236274 355807 236330 355816
rect 236012 354646 236132 354674
rect 236104 291854 236132 354646
rect 236092 291848 236144 291854
rect 236092 291790 236144 291796
rect 236288 279970 236316 355807
rect 237024 351898 237052 356215
rect 237012 351892 237064 351898
rect 237012 351834 237064 351840
rect 237010 351248 237066 351257
rect 237010 351183 237066 351192
rect 236644 341624 236696 341630
rect 236644 341566 236696 341572
rect 236656 279970 236684 341566
rect 237024 279970 237052 351183
rect 237378 348392 237434 348401
rect 237378 348327 237434 348336
rect 237392 279970 237420 348327
rect 238036 342242 238064 357167
rect 238758 357096 238814 357105
rect 238758 357031 238814 357040
rect 238116 355292 238168 355298
rect 238116 355234 238168 355240
rect 238024 342236 238076 342242
rect 238024 342178 238076 342184
rect 237748 341692 237800 341698
rect 237748 341634 237800 341640
rect 237760 279970 237788 341634
rect 238128 279970 238156 355234
rect 238772 352578 238800 357031
rect 239588 355292 239640 355298
rect 239588 355234 239640 355240
rect 238760 352572 238812 352578
rect 238760 352514 238812 352520
rect 238482 304192 238538 304201
rect 238482 304127 238538 304136
rect 238496 279970 238524 304127
rect 239220 293752 239272 293758
rect 239220 293694 239272 293700
rect 238852 290284 238904 290290
rect 238852 290226 238904 290232
rect 238864 279970 238892 290226
rect 239232 279970 239260 293694
rect 239600 279970 239628 355234
rect 239968 279970 239996 358430
rect 243636 358420 243688 358426
rect 243636 358362 243688 358368
rect 243542 357368 243598 357377
rect 243542 357303 243598 357312
rect 243556 356998 243584 357303
rect 243544 356992 243596 356998
rect 243544 356934 243596 356940
rect 240230 356008 240286 356017
rect 240230 355943 240286 355952
rect 240244 287978 240272 355943
rect 240322 355736 240378 355745
rect 240322 355671 240378 355680
rect 240232 287972 240284 287978
rect 240232 287914 240284 287920
rect 240336 279970 240364 355671
rect 241060 351212 241112 351218
rect 241060 351154 241112 351160
rect 240692 336048 240744 336054
rect 240692 335990 240744 335996
rect 240704 279970 240732 335990
rect 241072 279970 241100 351154
rect 241428 348492 241480 348498
rect 241428 348434 241480 348440
rect 241440 279970 241468 348434
rect 243556 345030 243584 356934
rect 243544 345024 243596 345030
rect 243544 344966 243596 344972
rect 243268 307080 243320 307086
rect 243268 307022 243320 307028
rect 242900 293684 242952 293690
rect 242900 293626 242952 293632
rect 242532 290352 242584 290358
rect 242532 290294 242584 290300
rect 242164 289196 242216 289202
rect 242164 289138 242216 289144
rect 241796 287904 241848 287910
rect 241796 287846 241848 287852
rect 241808 279970 241836 287846
rect 242176 279970 242204 289138
rect 242544 279970 242572 290294
rect 242912 279970 242940 293626
rect 243280 279970 243308 307022
rect 243648 279970 243676 358362
rect 246948 358352 247000 358358
rect 246948 358294 247000 358300
rect 244922 356960 244978 356969
rect 244922 356895 244978 356904
rect 245106 356960 245162 356969
rect 245106 356895 245162 356904
rect 244936 356658 244964 356895
rect 244924 356652 244976 356658
rect 244924 356594 244976 356600
rect 244280 356312 244332 356318
rect 244280 356254 244332 356260
rect 244292 355638 244320 356254
rect 244280 355632 244332 355638
rect 244002 355600 244058 355609
rect 244280 355574 244332 355580
rect 244002 355535 244058 355544
rect 244016 279970 244044 355535
rect 244292 286550 244320 355574
rect 244740 351280 244792 351286
rect 244740 351222 244792 351228
rect 244372 344412 244424 344418
rect 244372 344354 244424 344360
rect 244280 286544 244332 286550
rect 244280 286486 244332 286492
rect 244384 279970 244412 344354
rect 244752 279970 244780 351222
rect 244936 340882 244964 356594
rect 245120 356153 245148 356895
rect 245566 356688 245622 356697
rect 245566 356623 245622 356632
rect 245580 356318 245608 356623
rect 246854 356416 246910 356425
rect 246854 356351 246910 356360
rect 245568 356312 245620 356318
rect 245568 356254 245620 356260
rect 246868 356250 246896 356351
rect 245660 356244 245712 356250
rect 245660 356186 245712 356192
rect 246856 356244 246908 356250
rect 246856 356186 246908 356192
rect 245106 356144 245162 356153
rect 245106 356079 245162 356088
rect 245672 351354 245700 356186
rect 245660 351348 245712 351354
rect 245660 351290 245712 351296
rect 245108 348560 245160 348566
rect 245108 348502 245160 348508
rect 244924 340876 244976 340882
rect 244924 340818 244976 340824
rect 245120 279970 245148 348502
rect 245476 315444 245528 315450
rect 245476 315386 245528 315392
rect 245488 279970 245516 315386
rect 246212 293276 246264 293282
rect 246212 293218 246264 293224
rect 245844 290420 245896 290426
rect 245844 290362 245896 290368
rect 245856 279970 245884 290362
rect 246224 279970 246252 293218
rect 246580 291848 246632 291854
rect 246580 291790 246632 291796
rect 246592 279970 246620 291790
rect 246960 279970 246988 358294
rect 250260 358284 250312 358290
rect 250260 358226 250312 358232
rect 247222 357368 247278 357377
rect 247222 357303 247278 357312
rect 248694 357368 248750 357377
rect 248694 357303 248750 357312
rect 249982 357368 250038 357377
rect 249982 357303 250038 357312
rect 247130 356552 247186 356561
rect 247130 356487 247186 356496
rect 247144 356114 247172 356487
rect 247132 356108 247184 356114
rect 247132 356050 247184 356056
rect 247144 355366 247172 356050
rect 247132 355360 247184 355366
rect 247132 355302 247184 355308
rect 247144 285258 247172 355302
rect 247236 315382 247264 357303
rect 248708 356182 248736 357303
rect 249708 356788 249760 356794
rect 249708 356730 249760 356736
rect 249720 356182 249748 356730
rect 248696 356176 248748 356182
rect 248696 356118 248748 356124
rect 249708 356176 249760 356182
rect 249708 356118 249760 356124
rect 247314 355464 247370 355473
rect 247314 355399 247370 355408
rect 247224 315376 247276 315382
rect 247224 315318 247276 315324
rect 247132 285252 247184 285258
rect 247132 285194 247184 285200
rect 247328 279970 247356 355399
rect 248052 351348 248104 351354
rect 248052 351290 248104 351296
rect 247684 349852 247736 349858
rect 247684 349794 247736 349800
rect 247696 279970 247724 349794
rect 248064 279970 248092 351290
rect 248788 350532 248840 350538
rect 248788 350474 248840 350480
rect 248420 348628 248472 348634
rect 248420 348570 248472 348576
rect 248432 279970 248460 348570
rect 248800 279970 248828 350474
rect 249996 327894 250024 357303
rect 250074 356688 250130 356697
rect 250074 356623 250130 356632
rect 250088 356590 250116 356623
rect 250076 356584 250128 356590
rect 250076 356526 250128 356532
rect 250088 355502 250116 356526
rect 250076 355496 250128 355502
rect 250076 355438 250128 355444
rect 250088 341698 250116 355438
rect 250076 341692 250128 341698
rect 250076 341634 250128 341640
rect 249984 327888 250036 327894
rect 249984 327830 250036 327836
rect 249892 295996 249944 296002
rect 249892 295938 249944 295944
rect 249522 293584 249578 293593
rect 249522 293519 249578 293528
rect 248970 282568 249026 282577
rect 248970 282503 249026 282512
rect 248984 279970 249012 282503
rect 249536 279970 249564 293519
rect 249904 279970 249932 295938
rect 250272 279970 250300 358226
rect 253572 358216 253624 358222
rect 250626 358184 250682 358193
rect 253572 358158 253624 358164
rect 250626 358119 250682 358128
rect 250640 279970 250668 358119
rect 251270 357368 251326 357377
rect 251270 357303 251326 357312
rect 252650 357368 252706 357377
rect 252650 357303 252706 357312
rect 251284 356862 251312 357303
rect 251272 356856 251324 356862
rect 251272 356798 251324 356804
rect 251284 355570 251312 356798
rect 252100 356720 252152 356726
rect 252100 356662 252152 356668
rect 252282 356688 252338 356697
rect 251456 356380 251508 356386
rect 251456 356322 251508 356328
rect 251468 355842 251496 356322
rect 251456 355836 251508 355842
rect 251456 355778 251508 355784
rect 251272 355564 251324 355570
rect 251272 355506 251324 355512
rect 251088 355428 251140 355434
rect 251088 355370 251140 355376
rect 251100 354754 251128 355370
rect 251088 354748 251140 354754
rect 251088 354690 251140 354696
rect 251100 350538 251128 354690
rect 251088 350532 251140 350538
rect 251088 350474 251140 350480
rect 250996 337408 251048 337414
rect 250996 337350 251048 337356
rect 251008 279970 251036 337350
rect 251284 287910 251312 355506
rect 251362 354104 251418 354113
rect 251362 354039 251418 354048
rect 251272 287904 251324 287910
rect 251272 287846 251324 287852
rect 251376 279970 251404 354039
rect 251468 315450 251496 355778
rect 252112 353258 252140 356662
rect 252282 356623 252338 356632
rect 252296 356386 252324 356623
rect 252284 356380 252336 356386
rect 252284 356322 252336 356328
rect 252100 353252 252152 353258
rect 252100 353194 252152 353200
rect 251732 351416 251784 351422
rect 251732 351358 251784 351364
rect 251456 315444 251508 315450
rect 251456 315386 251508 315392
rect 251744 279970 251772 351358
rect 252112 279970 252140 353194
rect 252664 293826 252692 357303
rect 253386 356552 253442 356561
rect 253386 356487 253442 356496
rect 253400 356182 253428 356487
rect 252836 356176 252888 356182
rect 252836 356118 252888 356124
rect 253388 356176 253440 356182
rect 253388 356118 253440 356124
rect 252848 354754 252876 356118
rect 252836 354748 252888 354754
rect 252836 354690 252888 354696
rect 253204 351824 253256 351830
rect 253204 351766 253256 351772
rect 252652 293820 252704 293826
rect 252652 293762 252704 293768
rect 252834 290864 252890 290873
rect 252834 290799 252890 290808
rect 252284 282328 252336 282334
rect 252284 282270 252336 282276
rect 252296 279970 252324 282270
rect 252848 279970 252876 290799
rect 253216 279970 253244 351766
rect 253584 279970 253612 358158
rect 253938 358048 253994 358057
rect 253938 357983 253994 357992
rect 253952 279970 253980 357983
rect 254582 357368 254638 357377
rect 254582 357303 254638 357312
rect 255410 357368 255466 357377
rect 255410 357303 255466 357312
rect 254596 356726 254624 357303
rect 254584 356720 254636 356726
rect 254584 356662 254636 356668
rect 255320 356448 255372 356454
rect 255320 356390 255372 356396
rect 255332 355910 255360 356390
rect 255320 355904 255372 355910
rect 255320 355846 255372 355852
rect 255042 351384 255098 351393
rect 255042 351319 255098 351328
rect 254308 305652 254360 305658
rect 254308 305594 254360 305600
rect 254320 279970 254348 305594
rect 254676 297696 254728 297702
rect 254676 297638 254728 297644
rect 254688 279970 254716 297638
rect 255056 279970 255084 351319
rect 255332 279970 255360 355846
rect 255424 330682 255452 357303
rect 255778 356688 255834 356697
rect 255778 356623 255834 356632
rect 255792 356454 255820 356623
rect 255780 356448 255832 356454
rect 255780 356390 255832 356396
rect 255412 330676 255464 330682
rect 255412 330618 255464 330624
rect 256516 304428 256568 304434
rect 256516 304370 256568 304376
rect 256146 290728 256202 290737
rect 256146 290663 256202 290672
rect 255594 285424 255650 285433
rect 255594 285359 255650 285368
rect 255608 279970 255636 285359
rect 256160 279970 256188 290663
rect 256528 279970 256556 304370
rect 256896 279970 256924 359178
rect 257264 279970 257292 359246
rect 257342 357368 257398 357377
rect 257342 357303 257398 357312
rect 258170 357368 258226 357377
rect 258170 357303 258226 357312
rect 257356 356930 257384 357303
rect 257344 356924 257396 356930
rect 257344 356866 257396 356872
rect 257356 355706 257384 356866
rect 257344 355700 257396 355706
rect 257344 355642 257396 355648
rect 257356 342990 257384 355642
rect 257986 354240 258042 354249
rect 257986 354175 258042 354184
rect 257344 342984 257396 342990
rect 257344 342926 257396 342932
rect 257620 320952 257672 320958
rect 257620 320894 257672 320900
rect 257632 279970 257660 320894
rect 258000 279970 258028 354175
rect 258184 340270 258212 357303
rect 258814 356688 258870 356697
rect 258814 356623 258870 356632
rect 258828 356522 258856 356623
rect 258816 356516 258868 356522
rect 258816 356458 258868 356464
rect 258828 355774 258856 356458
rect 258816 355768 258868 355774
rect 258816 355710 258868 355716
rect 258828 354674 258856 355710
rect 258736 354646 258856 354674
rect 258264 342984 258316 342990
rect 258264 342926 258316 342932
rect 258172 340264 258224 340270
rect 258172 340206 258224 340212
rect 258276 282878 258304 342926
rect 258736 299470 258764 354646
rect 258724 299464 258776 299470
rect 258724 299406 258776 299412
rect 258356 298784 258408 298790
rect 258356 298726 258408 298732
rect 258264 282872 258316 282878
rect 258264 282814 258316 282820
rect 258368 279970 258396 298726
rect 259460 292052 259512 292058
rect 259460 291994 259512 292000
rect 258906 285288 258962 285297
rect 258906 285223 258962 285232
rect 258540 282872 258592 282878
rect 258540 282814 258592 282820
rect 258552 279970 258580 282814
rect 258920 279970 258948 285223
rect 259472 279970 259500 291994
rect 259748 282878 259776 359450
rect 260562 359272 260618 359281
rect 260562 359207 260618 359216
rect 260194 356688 260250 356697
rect 260194 356623 260250 356632
rect 260102 356416 260158 356425
rect 260102 356351 260158 356360
rect 260116 355978 260144 356351
rect 260208 356046 260236 356623
rect 260196 356040 260248 356046
rect 260196 355982 260248 355988
rect 260104 355972 260156 355978
rect 260104 355914 260156 355920
rect 259828 315376 259880 315382
rect 259828 315318 259880 315324
rect 259736 282872 259788 282878
rect 259736 282814 259788 282820
rect 259840 279970 259868 315318
rect 260116 285190 260144 355914
rect 260208 298110 260236 355982
rect 260196 298104 260248 298110
rect 260196 298046 260248 298052
rect 260104 285184 260156 285190
rect 260104 285126 260156 285132
rect 260012 282872 260064 282878
rect 260012 282814 260064 282820
rect 260024 279970 260052 282814
rect 260576 279970 260604 359207
rect 260838 357368 260894 357377
rect 260838 357303 260894 357312
rect 260852 354006 260880 357303
rect 260840 354000 260892 354006
rect 260840 353942 260892 353948
rect 260932 304292 260984 304298
rect 260932 304234 260984 304240
rect 260944 279970 260972 304234
rect 261312 279970 261340 359450
rect 262128 357400 262180 357406
rect 262126 357368 262128 357377
rect 262180 357368 262182 357377
rect 262126 357303 262182 357312
rect 262770 357368 262826 357377
rect 262770 357303 262772 357312
rect 262140 356998 262168 357303
rect 262824 357303 262826 357312
rect 262772 357274 262824 357280
rect 262128 356992 262180 356998
rect 262128 356934 262180 356940
rect 262784 356658 262812 357274
rect 262772 356652 262824 356658
rect 262772 356594 262824 356600
rect 261668 351484 261720 351490
rect 261668 351426 261720 351432
rect 261680 279970 261708 351426
rect 262036 299464 262088 299470
rect 262036 299406 262088 299412
rect 262048 279970 262076 299406
rect 263140 297492 263192 297498
rect 263140 297434 263192 297440
rect 262770 289096 262826 289105
rect 262770 289031 262826 289040
rect 262218 285152 262274 285161
rect 262218 285087 262274 285096
rect 262232 279970 262260 285087
rect 262784 279970 262812 289031
rect 263152 279970 263180 297434
rect 263520 279970 263548 359518
rect 263690 357368 263746 357377
rect 263690 357303 263746 357312
rect 263600 357264 263652 357270
rect 263600 357206 263652 357212
rect 263612 356318 263640 357206
rect 263600 356312 263652 356318
rect 263600 356254 263652 356260
rect 263704 304366 263732 357303
rect 263692 304360 263744 304366
rect 263692 304302 263744 304308
rect 263888 279970 263916 359615
rect 270132 359586 270184 359592
rect 264612 359576 264664 359582
rect 264612 359518 264664 359524
rect 263966 357368 264022 357377
rect 263966 357303 264022 357312
rect 263980 357270 264008 357303
rect 263968 357264 264020 357270
rect 263968 357206 264020 357212
rect 264244 293276 264296 293282
rect 264244 293218 264296 293224
rect 264256 279970 264284 293218
rect 264624 279970 264652 359518
rect 266634 359408 266690 359417
rect 266634 359343 266690 359352
rect 266820 359372 266872 359378
rect 265714 357368 265770 357377
rect 265714 357303 265770 357312
rect 266450 357368 266506 357377
rect 266450 357303 266506 357312
rect 265728 356998 265756 357303
rect 266360 357060 266412 357066
rect 266360 357002 266412 357008
rect 265072 356992 265124 356998
rect 265072 356934 265124 356940
rect 265716 356992 265768 356998
rect 265716 356934 265768 356940
rect 264978 356552 265034 356561
rect 264978 356487 265034 356496
rect 264992 355298 265020 356487
rect 265084 356250 265112 356934
rect 266372 356794 266400 357002
rect 266464 356794 266492 357303
rect 266360 356788 266412 356794
rect 266360 356730 266412 356736
rect 266452 356788 266504 356794
rect 266452 356730 266504 356736
rect 265072 356244 265124 356250
rect 265072 356186 265124 356192
rect 266464 356114 266492 356730
rect 266452 356108 266504 356114
rect 266452 356050 266504 356056
rect 264980 355292 265032 355298
rect 264980 355234 265032 355240
rect 264980 351552 265032 351558
rect 264980 351494 265032 351500
rect 264992 279970 265020 351494
rect 265348 298104 265400 298110
rect 265348 298046 265400 298052
rect 265360 279970 265388 298046
rect 266084 293616 266136 293622
rect 266084 293558 266136 293564
rect 265530 285016 265586 285025
rect 265530 284951 265586 284960
rect 265544 279970 265572 284951
rect 266096 279970 266124 293558
rect 266452 292052 266504 292058
rect 266452 291994 266504 292000
rect 266464 279970 266492 291994
rect 266648 282878 266676 359343
rect 266820 359314 266872 359320
rect 266636 282872 266688 282878
rect 266636 282814 266688 282820
rect 266832 279970 266860 359314
rect 267554 357368 267610 357377
rect 267554 357303 267610 357312
rect 267738 357368 267794 357377
rect 267738 357303 267794 357312
rect 268566 357368 268622 357377
rect 268566 357303 268622 357312
rect 269762 357368 269818 357377
rect 269762 357303 269818 357312
rect 267568 357066 267596 357303
rect 267556 357060 267608 357066
rect 267556 357002 267608 357008
rect 267556 316736 267608 316742
rect 267556 316678 267608 316684
rect 267004 282872 267056 282878
rect 267004 282814 267056 282820
rect 267016 279970 267044 282814
rect 267568 279970 267596 316678
rect 267752 307086 267780 357303
rect 268580 357202 268608 357303
rect 268292 357196 268344 357202
rect 268292 357138 268344 357144
rect 268568 357196 268620 357202
rect 268568 357138 268620 357144
rect 268304 356590 268332 357138
rect 269776 356862 269804 357303
rect 269764 356856 269816 356862
rect 269764 356798 269816 356804
rect 268292 356584 268344 356590
rect 268292 356526 268344 356532
rect 267922 354376 267978 354385
rect 267922 354311 267978 354320
rect 267740 307080 267792 307086
rect 267740 307022 267792 307028
rect 267936 279970 267964 354311
rect 269764 354204 269816 354210
rect 269764 354146 269816 354152
rect 268292 351620 268344 351626
rect 268292 351562 268344 351568
rect 268304 279970 268332 351562
rect 269396 291984 269448 291990
rect 269396 291926 269448 291932
rect 269026 287872 269082 287881
rect 269026 287807 269082 287816
rect 268476 285184 268528 285190
rect 268476 285126 268528 285132
rect 268488 279970 268516 285126
rect 269040 279970 269068 287807
rect 269408 279970 269436 291926
rect 269776 279970 269804 354146
rect 270144 279970 270172 359586
rect 270408 356856 270460 356862
rect 270408 356798 270460 356804
rect 270420 356318 270448 356798
rect 270408 356312 270460 356318
rect 270408 356254 270460 356260
rect 270512 279970 270540 359858
rect 273444 359848 273496 359854
rect 273444 359790 273496 359796
rect 279332 359848 279384 359854
rect 279332 359790 279384 359796
rect 273076 359712 273128 359718
rect 273076 359654 273128 359660
rect 271236 359644 271288 359650
rect 271236 359586 271288 359592
rect 270590 357368 270646 357377
rect 270590 357303 270646 357312
rect 271142 357368 271198 357377
rect 271142 357303 271198 357312
rect 270604 291854 270632 357303
rect 271156 356386 271184 357303
rect 271144 356380 271196 356386
rect 271144 356322 271196 356328
rect 270868 318096 270920 318102
rect 270868 318038 270920 318044
rect 270592 291848 270644 291854
rect 270592 291790 270644 291796
rect 270880 279970 270908 318038
rect 271248 279970 271276 359586
rect 272154 357368 272210 357377
rect 272154 357303 272210 357312
rect 272168 356862 272196 357303
rect 272156 356856 272208 356862
rect 272156 356798 272208 356804
rect 272168 356182 272196 356798
rect 272156 356176 272208 356182
rect 272156 356118 272208 356124
rect 271604 351688 271656 351694
rect 271604 351630 271656 351636
rect 271616 279970 271644 351630
rect 272340 295112 272392 295118
rect 272340 295054 272392 295060
rect 271970 287736 272026 287745
rect 271970 287671 272026 287680
rect 271984 279970 272012 287671
rect 272352 279970 272380 295054
rect 272708 293616 272760 293622
rect 272708 293558 272760 293564
rect 272720 279970 272748 293558
rect 273088 279970 273116 359654
rect 273350 357368 273406 357377
rect 273350 357303 273406 357312
rect 273364 356726 273392 357303
rect 273352 356720 273404 356726
rect 273352 356662 273404 356668
rect 273350 356144 273406 356153
rect 273350 356079 273406 356088
rect 273364 296002 273392 356079
rect 273352 295996 273404 296002
rect 273352 295938 273404 295944
rect 273456 279970 273484 359790
rect 276388 359780 276440 359786
rect 276388 359722 276440 359728
rect 276112 359440 276164 359446
rect 276112 359382 276164 359388
rect 276018 358184 276074 358193
rect 276018 358119 276074 358128
rect 274546 357368 274602 357377
rect 274546 357303 274602 357312
rect 275926 357368 275982 357377
rect 275926 357303 275982 357312
rect 274456 356720 274508 356726
rect 274456 356662 274508 356668
rect 274468 356250 274496 356662
rect 274560 356658 274588 357303
rect 275940 356930 275968 357303
rect 275928 356924 275980 356930
rect 275928 356866 275980 356872
rect 274548 356652 274600 356658
rect 274548 356594 274600 356600
rect 274560 356454 274588 356594
rect 275940 356590 275968 356866
rect 275928 356584 275980 356590
rect 275928 356526 275980 356532
rect 274548 356448 274600 356454
rect 274548 356390 274600 356396
rect 274456 356244 274508 356250
rect 274456 356186 274508 356192
rect 275652 355632 275704 355638
rect 275652 355574 275704 355580
rect 274178 354512 274234 354521
rect 274178 354447 274234 354456
rect 273812 300144 273864 300150
rect 273812 300086 273864 300092
rect 273824 279970 273852 300086
rect 274192 279970 274220 354447
rect 274548 351756 274600 351762
rect 274548 351698 274600 351704
rect 274560 279970 274588 351698
rect 275284 294976 275336 294982
rect 275284 294918 275336 294924
rect 274916 287836 274968 287842
rect 274916 287778 274968 287784
rect 274928 279970 274956 287778
rect 275296 279970 275324 294918
rect 275664 279970 275692 355574
rect 276032 351830 276060 358119
rect 276020 351824 276072 351830
rect 276020 351766 276072 351772
rect 276124 350534 276152 359382
rect 276032 350506 276152 350534
rect 276032 279970 276060 350506
rect 276400 279970 276428 359722
rect 277124 359712 277176 359718
rect 277124 359654 277176 359660
rect 277030 357368 277086 357377
rect 277030 357303 277086 357312
rect 277044 356522 277072 357303
rect 277032 356516 277084 356522
rect 277032 356458 277084 356464
rect 276756 301504 276808 301510
rect 276756 301446 276808 301452
rect 276768 279970 276796 301446
rect 277136 279970 277164 359654
rect 277398 356144 277454 356153
rect 277398 356079 277454 356088
rect 277412 304434 277440 356079
rect 278964 354680 279016 354686
rect 278964 354622 279016 354628
rect 277492 351824 277544 351830
rect 277492 351766 277544 351772
rect 277400 304428 277452 304434
rect 277400 304370 277452 304376
rect 277504 279970 277532 351766
rect 278596 304360 278648 304366
rect 278596 304302 278648 304308
rect 278228 294908 278280 294914
rect 278228 294850 278280 294856
rect 277860 287768 277912 287774
rect 277860 287710 277912 287716
rect 277872 279970 277900 287710
rect 278240 279970 278268 294850
rect 278608 279970 278636 304302
rect 278976 279970 279004 354622
rect 279344 279970 279372 359790
rect 300676 359780 300728 359786
rect 300676 359722 300728 359728
rect 285218 359544 285274 359553
rect 285218 359479 285274 359488
rect 282274 359408 282330 359417
rect 282274 359343 282330 359352
rect 280158 356144 280214 356153
rect 280158 356079 280214 356088
rect 280068 354000 280120 354006
rect 280068 353942 280120 353948
rect 279700 308440 279752 308446
rect 279700 308382 279752 308388
rect 279712 279970 279740 308382
rect 280080 279970 280108 353942
rect 280172 315382 280200 356079
rect 281908 355360 281960 355366
rect 281908 355302 281960 355308
rect 280436 351892 280488 351898
rect 280436 351834 280488 351840
rect 280160 315376 280212 315382
rect 280160 315318 280212 315324
rect 280448 279970 280476 351834
rect 281540 296132 281592 296138
rect 281540 296074 281592 296080
rect 281172 294772 281224 294778
rect 281172 294714 281224 294720
rect 280804 287700 280856 287706
rect 280804 287642 280856 287648
rect 280816 279970 280844 287642
rect 281184 279970 281212 294714
rect 281552 279970 281580 296074
rect 281920 279970 281948 355302
rect 282288 279970 282316 359343
rect 282918 357368 282974 357377
rect 282918 357303 282974 357312
rect 282644 307080 282696 307086
rect 282644 307022 282696 307028
rect 282656 279970 282684 307022
rect 282932 297498 282960 357303
rect 284852 355428 284904 355434
rect 284852 355370 284904 355376
rect 283012 354068 283064 354074
rect 283012 354010 283064 354016
rect 282920 297492 282972 297498
rect 282920 297434 282972 297440
rect 283024 279970 283052 354010
rect 283380 351144 283432 351150
rect 283380 351086 283432 351092
rect 283392 279970 283420 351086
rect 284484 329180 284536 329186
rect 284484 329122 284536 329128
rect 284116 294840 284168 294846
rect 284116 294782 284168 294788
rect 283748 291168 283800 291174
rect 283748 291110 283800 291116
rect 283760 279970 283788 291110
rect 284128 279970 284156 294782
rect 284496 279970 284524 329122
rect 284864 279970 284892 355370
rect 285232 279970 285260 359479
rect 299572 358352 299624 358358
rect 299572 358294 299624 358300
rect 299938 358320 299994 358329
rect 296628 358284 296680 358290
rect 296628 358226 296680 358232
rect 293684 358216 293736 358222
rect 293684 358158 293736 358164
rect 285678 357368 285734 357377
rect 285678 357303 285734 357312
rect 287058 357368 287114 357377
rect 287058 357303 287114 357312
rect 289910 357368 289966 357377
rect 289910 357303 289966 357312
rect 292578 357368 292634 357377
rect 292578 357303 292634 357312
rect 285588 315376 285640 315382
rect 285588 315318 285640 315324
rect 285600 279970 285628 315318
rect 285692 292058 285720 357303
rect 287072 354210 287100 357303
rect 287796 355496 287848 355502
rect 287796 355438 287848 355444
rect 287060 354204 287112 354210
rect 287060 354146 287112 354152
rect 285956 354136 286008 354142
rect 285956 354078 286008 354084
rect 285680 292052 285732 292058
rect 285680 291994 285732 292000
rect 285968 279970 285996 354078
rect 286324 348696 286376 348702
rect 286324 348638 286376 348644
rect 286336 279970 286364 348638
rect 287060 295044 287112 295050
rect 287060 294986 287112 294992
rect 286692 291100 286744 291106
rect 286692 291042 286744 291048
rect 286704 279970 286732 291042
rect 287072 279970 287100 294986
rect 287428 291984 287480 291990
rect 287428 291926 287480 291932
rect 287440 279970 287468 291926
rect 287808 279970 287836 355438
rect 288900 354204 288952 354210
rect 288900 354146 288952 354152
rect 288164 353932 288216 353938
rect 288164 353874 288216 353880
rect 288176 279970 288204 353874
rect 288532 302932 288584 302938
rect 288532 302874 288584 302880
rect 288544 279970 288572 302874
rect 288912 279970 288940 354146
rect 289268 348764 289320 348770
rect 289268 348706 289320 348712
rect 289280 279970 289308 348706
rect 289924 293622 289952 357303
rect 292592 355638 292620 357303
rect 292580 355632 292632 355638
rect 292580 355574 292632 355580
rect 290740 355564 290792 355570
rect 290740 355506 290792 355512
rect 290004 296268 290056 296274
rect 290004 296210 290056 296216
rect 289912 293616 289964 293622
rect 289912 293558 289964 293564
rect 289636 291032 289688 291038
rect 289636 290974 289688 290980
rect 289648 279970 289676 290974
rect 290016 279970 290044 296210
rect 290372 293616 290424 293622
rect 290372 293558 290424 293564
rect 290384 279970 290412 293558
rect 290752 279970 290780 355506
rect 291844 354272 291896 354278
rect 291844 354214 291896 354220
rect 291108 353864 291160 353870
rect 291108 353806 291160 353812
rect 291120 279970 291148 353806
rect 291476 291848 291528 291854
rect 291476 291790 291528 291796
rect 291488 279970 291516 291790
rect 291856 279970 291884 354214
rect 292212 348832 292264 348838
rect 292212 348774 292264 348780
rect 292224 279970 292252 348774
rect 292946 293448 293002 293457
rect 292946 293383 293002 293392
rect 292580 290964 292632 290970
rect 292580 290906 292632 290912
rect 292592 279970 292620 290906
rect 292960 279970 292988 293383
rect 293316 292052 293368 292058
rect 293316 291994 293368 292000
rect 293328 279970 293356 291994
rect 293696 279970 293724 358158
rect 294050 358048 294106 358057
rect 294050 357983 294106 357992
rect 294064 279970 294092 357983
rect 295338 357368 295394 357377
rect 295338 357303 295394 357312
rect 294788 354340 294840 354346
rect 294788 354282 294840 354288
rect 294420 297492 294472 297498
rect 294420 297434 294472 297440
rect 294432 279970 294460 297434
rect 294800 279970 294828 354282
rect 295156 348900 295208 348906
rect 295156 348842 295208 348848
rect 295168 279970 295196 348842
rect 295352 304366 295380 357303
rect 295340 304360 295392 304366
rect 295340 304302 295392 304308
rect 296260 294636 296312 294642
rect 296260 294578 296312 294584
rect 295892 293548 295944 293554
rect 295892 293490 295944 293496
rect 295524 290896 295576 290902
rect 295524 290838 295576 290844
rect 295536 279970 295564 290838
rect 295904 279970 295932 293490
rect 296272 279970 296300 294578
rect 296640 279970 296668 358226
rect 296994 357912 297050 357921
rect 296994 357847 297050 357856
rect 297008 279970 297036 357847
rect 298190 357368 298246 357377
rect 298190 357303 298246 357312
rect 297732 354408 297784 354414
rect 297732 354350 297784 354356
rect 297364 295996 297416 296002
rect 297364 295938 297416 295944
rect 297376 279970 297404 295938
rect 297744 279970 297772 354350
rect 298100 348968 298152 348974
rect 298100 348910 298152 348916
rect 298112 279970 298140 348910
rect 298204 296138 298232 357303
rect 298192 296132 298244 296138
rect 298192 296074 298244 296080
rect 299204 296132 299256 296138
rect 299204 296074 299256 296080
rect 298836 293480 298888 293486
rect 298836 293422 298888 293428
rect 298468 290828 298520 290834
rect 298468 290770 298520 290776
rect 298480 279970 298508 290770
rect 298848 279970 298876 293422
rect 299216 279970 299244 296074
rect 299584 279970 299612 358294
rect 299938 358255 299994 358264
rect 299952 279970 299980 358255
rect 300308 311160 300360 311166
rect 300308 311102 300360 311108
rect 300320 279970 300348 311102
rect 300688 279970 300716 359722
rect 308770 358592 308826 358601
rect 305460 358556 305512 358562
rect 308770 358527 308826 358536
rect 305460 358498 305512 358504
rect 302516 358488 302568 358494
rect 302516 358430 302568 358436
rect 300858 358184 300914 358193
rect 300858 358119 300914 358128
rect 301042 358184 301098 358193
rect 301042 358119 301098 358128
rect 300872 329186 300900 358119
rect 301056 357921 301084 358119
rect 301042 357912 301098 357921
rect 301042 357847 301098 357856
rect 302238 357368 302294 357377
rect 302238 357303 302294 357312
rect 301044 349036 301096 349042
rect 301044 348978 301096 348984
rect 300860 329180 300912 329186
rect 300860 329122 300912 329128
rect 301056 279970 301084 348978
rect 301780 293412 301832 293418
rect 301780 293354 301832 293360
rect 301412 290760 301464 290766
rect 301412 290702 301464 290708
rect 301424 279970 301452 290702
rect 301792 279970 301820 293354
rect 302148 292120 302200 292126
rect 302148 292062 302200 292068
rect 302160 279970 302188 292062
rect 302252 291990 302280 357303
rect 302240 291984 302292 291990
rect 302240 291926 302292 291932
rect 302528 279970 302556 358430
rect 302884 358420 302936 358426
rect 302884 358362 302936 358368
rect 302896 279970 302924 358362
rect 304998 357368 305054 357377
rect 304998 357303 305054 357312
rect 303620 354476 303672 354482
rect 303620 354418 303672 354424
rect 303252 309800 303304 309806
rect 303252 309742 303304 309748
rect 303264 279970 303292 309742
rect 303632 279970 303660 354418
rect 303988 349104 304040 349110
rect 303988 349046 304040 349052
rect 304000 279970 304028 349046
rect 304724 296200 304776 296206
rect 304724 296142 304776 296148
rect 304356 290692 304408 290698
rect 304356 290634 304408 290640
rect 304368 279970 304396 290634
rect 304736 279970 304764 296142
rect 305012 293622 305040 357303
rect 305092 297764 305144 297770
rect 305092 297706 305144 297712
rect 305000 293616 305052 293622
rect 305000 293558 305052 293564
rect 305104 279970 305132 297706
rect 305472 279970 305500 358498
rect 305826 358456 305882 358465
rect 305826 358391 305882 358400
rect 305840 279970 305868 358391
rect 308404 358012 308456 358018
rect 308404 357954 308456 357960
rect 307758 357368 307814 357377
rect 307758 357303 307814 357312
rect 306564 354544 306616 354550
rect 306564 354486 306616 354492
rect 306196 319524 306248 319530
rect 306196 319466 306248 319472
rect 306208 279970 306236 319466
rect 306576 279970 306604 354486
rect 306932 348356 306984 348362
rect 306932 348298 306984 348304
rect 306944 279970 306972 348298
rect 307668 293344 307720 293350
rect 307668 293286 307720 293292
rect 307300 290624 307352 290630
rect 307300 290566 307352 290572
rect 307312 279970 307340 290566
rect 307680 279970 307708 293286
rect 307772 292058 307800 357303
rect 308036 293344 308088 293350
rect 308036 293286 308088 293292
rect 307760 292052 307812 292058
rect 307760 291994 307812 292000
rect 308048 279970 308076 293286
rect 308416 279970 308444 357954
rect 308784 279970 308812 358527
rect 311348 357944 311400 357950
rect 311348 357886 311400 357892
rect 310518 357368 310574 357377
rect 310518 357303 310574 357312
rect 309508 354612 309560 354618
rect 309508 354554 309560 354560
rect 309140 313948 309192 313954
rect 309140 313890 309192 313896
rect 309152 279970 309180 313890
rect 309520 279970 309548 354554
rect 309876 348288 309928 348294
rect 309876 348230 309928 348236
rect 309888 279970 309916 348230
rect 310532 294642 310560 357303
rect 310980 355632 311032 355638
rect 310980 355574 311032 355580
rect 310612 296064 310664 296070
rect 310612 296006 310664 296012
rect 310520 294636 310572 294642
rect 310520 294578 310572 294584
rect 310244 290556 310296 290562
rect 310244 290498 310296 290504
rect 310256 279970 310284 290498
rect 310624 279970 310652 296006
rect 310992 279970 311020 355574
rect 311360 279970 311388 357886
rect 311728 279970 311756 359858
rect 314292 359440 314344 359446
rect 314292 359382 314344 359388
rect 313278 357368 313334 357377
rect 313278 357303 313334 357312
rect 312452 351076 312504 351082
rect 312452 351018 312504 351024
rect 312084 290488 312136 290494
rect 312084 290430 312136 290436
rect 312096 279970 312124 290430
rect 312464 279970 312492 351018
rect 312820 348220 312872 348226
rect 312820 348162 312872 348168
rect 312832 279970 312860 348162
rect 313292 296138 313320 357303
rect 313924 353796 313976 353802
rect 313924 353738 313976 353744
rect 313280 296132 313332 296138
rect 313280 296074 313332 296080
rect 313554 293312 313610 293321
rect 313554 293247 313610 293256
rect 313188 290216 313240 290222
rect 313188 290158 313240 290164
rect 313200 279970 313228 290158
rect 313568 279970 313596 293247
rect 313936 279970 313964 353738
rect 314304 279970 314332 359382
rect 325698 358728 325754 358737
rect 325698 358663 325754 358672
rect 314660 357876 314712 357882
rect 314660 357818 314712 357824
rect 314672 279970 314700 357818
rect 314750 357368 314806 357377
rect 314750 357303 314806 357312
rect 317418 357368 317474 357377
rect 317418 357303 317474 357312
rect 320178 357368 320234 357377
rect 320178 357303 320234 357312
rect 314764 292126 314792 357303
rect 315396 351008 315448 351014
rect 315396 350950 315448 350956
rect 315028 294636 315080 294642
rect 315028 294578 315080 294584
rect 314752 292120 314804 292126
rect 314752 292062 314804 292068
rect 314844 282056 314896 282062
rect 314844 281998 314896 282004
rect 230032 279942 230092 279970
rect 230400 279942 230460 279970
rect 230584 279942 230828 279970
rect 231136 279942 231196 279970
rect 231504 279942 231564 279970
rect 231872 279942 231932 279970
rect 232240 279942 232300 279970
rect 232608 279942 232668 279970
rect 232976 279942 233036 279970
rect 233344 279942 233404 279970
rect 233712 279942 233772 279970
rect 234080 279942 234140 279970
rect 234448 279942 234508 279970
rect 234816 279942 234876 279970
rect 235184 279942 235244 279970
rect 235552 279942 235612 279970
rect 235920 279942 235980 279970
rect 236288 279942 236348 279970
rect 236656 279942 236716 279970
rect 237024 279942 237084 279970
rect 237392 279942 237452 279970
rect 237760 279942 237820 279970
rect 238128 279942 238188 279970
rect 238496 279942 238556 279970
rect 238864 279942 238924 279970
rect 239232 279942 239292 279970
rect 239600 279942 239660 279970
rect 239968 279942 240028 279970
rect 240336 279942 240396 279970
rect 240704 279942 240764 279970
rect 241072 279942 241132 279970
rect 241440 279942 241500 279970
rect 241808 279942 241868 279970
rect 242176 279942 242236 279970
rect 242544 279942 242604 279970
rect 242912 279942 242972 279970
rect 243280 279942 243340 279970
rect 243648 279942 243708 279970
rect 244016 279942 244076 279970
rect 244384 279942 244444 279970
rect 244752 279942 244812 279970
rect 245120 279942 245180 279970
rect 245488 279942 245548 279970
rect 245856 279942 245916 279970
rect 246224 279942 246284 279970
rect 246592 279942 246652 279970
rect 246960 279942 247020 279970
rect 247328 279942 247388 279970
rect 247696 279942 247756 279970
rect 248064 279942 248124 279970
rect 248432 279942 248492 279970
rect 248800 279942 248860 279970
rect 248984 279942 249228 279970
rect 249536 279942 249596 279970
rect 249904 279942 249964 279970
rect 250272 279942 250332 279970
rect 250640 279942 250700 279970
rect 251008 279942 251068 279970
rect 251376 279942 251436 279970
rect 251744 279942 251804 279970
rect 252112 279942 252172 279970
rect 252296 279942 252540 279970
rect 252848 279942 252908 279970
rect 253216 279942 253276 279970
rect 253584 279942 253644 279970
rect 253952 279942 254012 279970
rect 254320 279942 254380 279970
rect 254688 279942 254748 279970
rect 255056 279942 255116 279970
rect 255332 279942 255484 279970
rect 255608 279942 255852 279970
rect 256160 279942 256220 279970
rect 256528 279942 256588 279970
rect 256896 279942 256956 279970
rect 257264 279942 257324 279970
rect 257632 279942 257692 279970
rect 258000 279942 258060 279970
rect 258368 279942 258428 279970
rect 258552 279942 258796 279970
rect 258920 279942 259164 279970
rect 259472 279942 259532 279970
rect 259840 279942 259900 279970
rect 260024 279942 260268 279970
rect 260576 279942 260636 279970
rect 260944 279942 261004 279970
rect 261312 279942 261372 279970
rect 261680 279942 261740 279970
rect 262048 279942 262108 279970
rect 262232 279942 262476 279970
rect 262784 279942 262844 279970
rect 263152 279942 263212 279970
rect 263520 279942 263580 279970
rect 263888 279942 263948 279970
rect 264256 279942 264316 279970
rect 264624 279942 264684 279970
rect 264992 279942 265052 279970
rect 265360 279942 265420 279970
rect 265544 279942 265788 279970
rect 266096 279942 266156 279970
rect 266464 279942 266524 279970
rect 266832 279942 266892 279970
rect 267016 279942 267260 279970
rect 267568 279942 267628 279970
rect 267936 279942 267996 279970
rect 268304 279942 268364 279970
rect 268488 279942 268732 279970
rect 269040 279942 269100 279970
rect 269408 279942 269468 279970
rect 269776 279942 269836 279970
rect 270144 279942 270204 279970
rect 270512 279942 270572 279970
rect 270880 279942 270940 279970
rect 271248 279942 271308 279970
rect 271616 279942 271676 279970
rect 271984 279942 272044 279970
rect 272352 279942 272412 279970
rect 272720 279942 272780 279970
rect 273088 279942 273148 279970
rect 273456 279942 273516 279970
rect 273824 279942 273884 279970
rect 274192 279942 274252 279970
rect 274560 279942 274620 279970
rect 274928 279942 274988 279970
rect 275296 279942 275356 279970
rect 275664 279942 275724 279970
rect 276032 279942 276092 279970
rect 276400 279942 276460 279970
rect 276768 279942 276828 279970
rect 277136 279942 277196 279970
rect 277504 279942 277564 279970
rect 277872 279942 277932 279970
rect 278240 279942 278300 279970
rect 278608 279942 278668 279970
rect 278976 279942 279036 279970
rect 279344 279942 279404 279970
rect 279712 279942 279772 279970
rect 280080 279942 280140 279970
rect 280448 279942 280508 279970
rect 280816 279942 280876 279970
rect 281184 279942 281244 279970
rect 281552 279942 281612 279970
rect 281920 279942 281980 279970
rect 282288 279942 282348 279970
rect 282656 279942 282716 279970
rect 283024 279942 283084 279970
rect 283392 279942 283452 279970
rect 283760 279942 283820 279970
rect 284128 279942 284188 279970
rect 284496 279942 284556 279970
rect 284864 279942 284924 279970
rect 285232 279942 285292 279970
rect 285600 279942 285660 279970
rect 285968 279942 286028 279970
rect 286336 279942 286396 279970
rect 286704 279942 286764 279970
rect 287072 279942 287132 279970
rect 287440 279942 287500 279970
rect 287808 279942 287868 279970
rect 288176 279942 288236 279970
rect 288544 279942 288604 279970
rect 288912 279942 288972 279970
rect 289280 279942 289340 279970
rect 289648 279942 289708 279970
rect 290016 279942 290076 279970
rect 290384 279942 290444 279970
rect 290752 279942 290812 279970
rect 291120 279942 291180 279970
rect 291488 279942 291548 279970
rect 291856 279942 291916 279970
rect 292224 279942 292284 279970
rect 292592 279942 292652 279970
rect 292960 279942 293020 279970
rect 293328 279942 293388 279970
rect 293696 279942 293756 279970
rect 294064 279942 294124 279970
rect 294432 279942 294492 279970
rect 294800 279942 294860 279970
rect 295168 279942 295228 279970
rect 295536 279942 295596 279970
rect 295904 279942 295964 279970
rect 296272 279942 296332 279970
rect 296640 279942 296700 279970
rect 297008 279942 297068 279970
rect 297376 279942 297436 279970
rect 297744 279942 297804 279970
rect 298112 279942 298172 279970
rect 298480 279942 298540 279970
rect 298848 279942 298908 279970
rect 299216 279942 299276 279970
rect 299584 279942 299644 279970
rect 299952 279942 300012 279970
rect 300320 279942 300380 279970
rect 300688 279942 300748 279970
rect 301056 279942 301116 279970
rect 301424 279942 301484 279970
rect 301792 279942 301852 279970
rect 302160 279942 302220 279970
rect 302528 279942 302588 279970
rect 302896 279942 302956 279970
rect 303264 279942 303324 279970
rect 303632 279942 303692 279970
rect 304000 279942 304060 279970
rect 304368 279942 304428 279970
rect 304736 279942 304796 279970
rect 305104 279942 305164 279970
rect 305472 279942 305532 279970
rect 305840 279942 305900 279970
rect 306208 279942 306268 279970
rect 306576 279942 306636 279970
rect 306944 279942 307004 279970
rect 307312 279942 307372 279970
rect 307680 279942 307740 279970
rect 308048 279942 308108 279970
rect 308416 279942 308476 279970
rect 308784 279942 308844 279970
rect 309152 279942 309212 279970
rect 309520 279942 309580 279970
rect 309888 279942 309948 279970
rect 310256 279942 310316 279970
rect 310624 279942 310684 279970
rect 310992 279942 311052 279970
rect 311360 279942 311420 279970
rect 311728 279942 311788 279970
rect 312096 279942 312156 279970
rect 312464 279942 312524 279970
rect 312832 279942 312892 279970
rect 313200 279942 313260 279970
rect 313568 279942 313628 279970
rect 313936 279942 313996 279970
rect 314304 279942 314364 279970
rect 314672 279942 314732 279970
rect 314856 279886 314884 281998
rect 315040 279970 315068 294578
rect 315408 279970 315436 350950
rect 316682 342952 316738 342961
rect 316682 342887 316738 342896
rect 316696 289814 316724 342887
rect 317432 297770 317460 357303
rect 317420 297764 317472 297770
rect 317420 297706 317472 297712
rect 320192 293350 320220 357303
rect 322938 356144 322994 356153
rect 322938 356079 322994 356088
rect 322952 355638 322980 356079
rect 322940 355632 322992 355638
rect 322940 355574 322992 355580
rect 325712 353802 325740 358663
rect 356624 358057 356652 596362
rect 356702 476776 356758 476785
rect 356702 476711 356758 476720
rect 356610 358048 356666 358057
rect 356610 357983 356666 357992
rect 325700 353796 325752 353802
rect 325700 353738 325752 353744
rect 356716 297702 356744 476711
rect 356808 298790 356836 596799
rect 357900 596770 357952 596776
rect 357716 596692 357768 596698
rect 357716 596634 357768 596640
rect 357532 596624 357584 596630
rect 357532 596566 357584 596572
rect 357440 596352 357492 596358
rect 357440 596294 357492 596300
rect 356886 477048 356942 477057
rect 356886 476983 356942 476992
rect 356796 298784 356848 298790
rect 356796 298726 356848 298732
rect 356704 297696 356756 297702
rect 356704 297638 356756 297644
rect 356900 297566 356928 476983
rect 357070 476912 357126 476921
rect 356980 476876 357032 476882
rect 357070 476847 357126 476856
rect 356980 476818 357032 476824
rect 356992 357950 357020 476818
rect 356980 357944 357032 357950
rect 356980 357886 357032 357892
rect 357084 297634 357112 476847
rect 357164 476468 357216 476474
rect 357164 476410 357216 476416
rect 357176 358222 357204 476410
rect 357164 358216 357216 358222
rect 357164 358158 357216 358164
rect 357452 353870 357480 596294
rect 357544 358329 357572 596566
rect 357624 596488 357676 596494
rect 357624 596430 357676 596436
rect 357530 358320 357586 358329
rect 357530 358255 357586 358264
rect 357636 358193 357664 596430
rect 357728 358465 357756 596634
rect 357808 596216 357860 596222
rect 357808 596158 357860 596164
rect 357820 359854 357848 596158
rect 357912 359922 357940 596770
rect 358832 560289 358860 678943
rect 359004 596896 359056 596902
rect 359004 596838 359056 596844
rect 358912 596284 358964 596290
rect 358912 596226 358964 596232
rect 358818 560280 358874 560289
rect 358818 560215 358874 560224
rect 358176 476672 358228 476678
rect 358176 476614 358228 476620
rect 358084 476536 358136 476542
rect 358084 476478 358136 476484
rect 357992 476128 358044 476134
rect 357992 476070 358044 476076
rect 357900 359916 357952 359922
rect 357900 359858 357952 359864
rect 357808 359848 357860 359854
rect 357808 359790 357860 359796
rect 357714 358456 357770 358465
rect 357714 358391 357770 358400
rect 357622 358184 357678 358193
rect 357622 358119 357678 358128
rect 358004 354686 358032 476070
rect 358096 358290 358124 476478
rect 358188 358494 358216 476614
rect 358820 454776 358872 454782
rect 358820 454718 358872 454724
rect 358832 453354 358860 454718
rect 358820 453348 358872 453354
rect 358820 453290 358872 453296
rect 358832 439249 358860 453290
rect 358818 439240 358874 439249
rect 358818 439175 358874 439184
rect 358268 367124 358320 367130
rect 358268 367066 358320 367072
rect 358176 358488 358228 358494
rect 358176 358430 358228 358436
rect 358084 358284 358136 358290
rect 358084 358226 358136 358232
rect 357992 354680 358044 354686
rect 357992 354622 358044 354628
rect 357440 353864 357492 353870
rect 357440 353806 357492 353812
rect 357072 297628 357124 297634
rect 357072 297570 357124 297576
rect 356888 297560 356940 297566
rect 356888 297502 356940 297508
rect 320180 293344 320232 293350
rect 320180 293286 320232 293292
rect 358280 291922 358308 367066
rect 358268 291916 358320 291922
rect 358268 291858 358320 291864
rect 316684 289808 316736 289814
rect 316684 289750 316736 289756
rect 316696 289066 316724 289750
rect 316132 289060 316184 289066
rect 316132 289002 316184 289008
rect 316684 289060 316736 289066
rect 316684 289002 316736 289008
rect 315762 282296 315818 282305
rect 315762 282231 315818 282240
rect 315776 279970 315804 282231
rect 316144 279970 316172 289002
rect 319536 287632 319588 287638
rect 319536 287574 319588 287580
rect 318156 282124 318208 282130
rect 318156 282066 318208 282072
rect 318064 281104 318116 281110
rect 318064 281046 318116 281052
rect 315040 279942 315100 279970
rect 315408 279942 315468 279970
rect 315776 279942 315836 279970
rect 316144 279942 316204 279970
rect 314844 279880 314896 279886
rect 211632 279806 211692 279834
rect 314844 279822 314896 279828
rect 187884 279744 187936 279750
rect 177468 279682 177712 279698
rect 187884 279686 187936 279692
rect 177468 279676 177724 279682
rect 177468 279670 177672 279676
rect 177672 279618 177724 279624
rect 158812 279608 158864 279614
rect 123850 279576 123906 279585
rect 123906 279534 124108 279562
rect 180616 279608 180668 279614
rect 158812 279550 158864 279556
rect 180412 279556 180616 279562
rect 183928 279608 183980 279614
rect 180412 279550 180668 279556
rect 183724 279556 183928 279562
rect 183724 279550 183980 279556
rect 180412 279534 180656 279550
rect 183724 279534 183968 279550
rect 123850 279511 123906 279520
rect 123712 279304 123768 279313
rect 123712 279239 123768 279248
rect 318076 232529 318104 281046
rect 318168 233889 318196 282066
rect 319444 281988 319496 281994
rect 319444 281930 319496 281936
rect 318248 281036 318300 281042
rect 318248 280978 318300 280984
rect 318260 271969 318288 280978
rect 318246 271960 318302 271969
rect 318246 271895 318302 271904
rect 319456 233918 319484 281930
rect 319444 233912 319496 233918
rect 318154 233880 318210 233889
rect 319444 233854 319496 233860
rect 318154 233815 318210 233824
rect 319548 232762 319576 287574
rect 319720 287564 319772 287570
rect 319720 287506 319772 287512
rect 319626 287464 319682 287473
rect 319626 287399 319682 287408
rect 319536 232756 319588 232762
rect 319536 232698 319588 232704
rect 319640 232558 319668 287399
rect 319732 232830 319760 287506
rect 320822 287328 320878 287337
rect 320822 287263 320878 287272
rect 319904 282260 319956 282266
rect 319904 282202 319956 282208
rect 319810 282160 319866 282169
rect 319810 282095 319866 282104
rect 319720 232824 319772 232830
rect 319720 232766 319772 232772
rect 319824 232626 319852 282095
rect 319916 232898 319944 282202
rect 320088 282192 320140 282198
rect 320088 282134 320140 282140
rect 319996 280696 320048 280702
rect 319996 280638 320048 280644
rect 320008 233238 320036 280638
rect 320100 233986 320128 282134
rect 320088 233980 320140 233986
rect 320088 233922 320140 233928
rect 319996 233232 320048 233238
rect 319996 233174 320048 233180
rect 319904 232892 319956 232898
rect 319904 232834 319956 232840
rect 320836 232694 320864 287263
rect 321100 283824 321152 283830
rect 321100 283766 321152 283772
rect 320916 281920 320968 281926
rect 320916 281862 320968 281868
rect 320928 232966 320956 281862
rect 321008 281852 321060 281858
rect 321008 281794 321060 281800
rect 321020 233034 321048 281794
rect 321112 245614 321140 283766
rect 321192 280764 321244 280770
rect 321192 280706 321244 280712
rect 321204 259418 321232 280706
rect 321192 259412 321244 259418
rect 321192 259354 321244 259360
rect 321100 245608 321152 245614
rect 321100 245550 321152 245556
rect 321008 233028 321060 233034
rect 321008 232970 321060 232976
rect 320916 232960 320968 232966
rect 320916 232902 320968 232908
rect 320824 232688 320876 232694
rect 320824 232630 320876 232636
rect 319812 232620 319864 232626
rect 319812 232562 319864 232568
rect 319628 232552 319680 232558
rect 318062 232520 318118 232529
rect 319628 232494 319680 232500
rect 318062 232455 318118 232464
rect 319444 231872 319496 231878
rect 319444 231814 319496 231820
rect 318062 230616 318118 230625
rect 318062 230551 318118 230560
rect 318076 80646 318104 230551
rect 318154 229120 318210 229129
rect 318154 229055 318210 229064
rect 318168 93854 318196 229055
rect 318168 93826 318380 93854
rect 314108 80640 314160 80646
rect 313812 80588 314108 80594
rect 313812 80582 314160 80588
rect 318064 80640 318116 80646
rect 318064 80582 318116 80588
rect 313812 80566 314148 80582
rect 121656 80022 121992 80050
rect 123036 80022 123372 80050
rect 124752 80022 125088 80050
rect 121656 77994 121684 80022
rect 123036 78062 123064 80022
rect 123024 78056 123076 78062
rect 123024 77998 123076 78004
rect 121644 77988 121696 77994
rect 121644 77930 121696 77936
rect 125060 77314 125088 80022
rect 125704 80022 126132 80050
rect 127084 80022 127512 80050
rect 128892 80022 129228 80050
rect 125048 77308 125100 77314
rect 125048 77250 125100 77256
rect 125600 77308 125652 77314
rect 125600 77250 125652 77256
rect 121368 20664 121420 20670
rect 121368 20606 121420 20612
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 120724 6860 120776 6866
rect 120724 6802 120776 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 77250
rect 125704 3466 125732 80022
rect 127084 6914 127112 80022
rect 129200 77314 129228 80022
rect 129844 80022 130272 80050
rect 131132 80022 131652 80050
rect 132512 80022 133032 80050
rect 133984 80022 134412 80050
rect 135272 80022 135792 80050
rect 136652 80022 137172 80050
rect 138032 80022 138552 80050
rect 139412 80022 139932 80050
rect 140792 80022 141312 80050
rect 142172 80022 142692 80050
rect 143552 80022 144072 80050
rect 144932 80022 145452 80050
rect 146312 80022 146832 80050
rect 147692 80022 148212 80050
rect 149072 80022 149592 80050
rect 150452 80022 150972 80050
rect 151832 80022 152352 80050
rect 153212 80022 153732 80050
rect 155112 80022 155448 80050
rect 156492 80022 156828 80050
rect 157872 80022 158208 80050
rect 159252 80022 159588 80050
rect 160632 80022 160968 80050
rect 162012 80022 162348 80050
rect 163392 80022 163728 80050
rect 164772 80022 165108 80050
rect 129188 77308 129240 77314
rect 129188 77250 129240 77256
rect 129740 77308 129792 77314
rect 129740 77250 129792 77256
rect 126992 6886 127112 6914
rect 125692 3460 125744 3466
rect 125692 3402 125744 3408
rect 126992 480 127020 6886
rect 129752 3482 129780 77250
rect 129844 4146 129872 80022
rect 129832 4140 129884 4146
rect 129832 4082 129884 4088
rect 131132 3670 131160 80022
rect 131120 3664 131172 3670
rect 131120 3606 131172 3612
rect 128176 3460 128228 3466
rect 129752 3454 130608 3482
rect 132512 3466 132540 80022
rect 133984 3602 134012 80022
rect 134156 4140 134208 4146
rect 134156 4082 134208 4088
rect 133972 3596 134024 3602
rect 133972 3538 134024 3544
rect 128176 3402 128228 3408
rect 128188 480 128216 3402
rect 130580 480 130608 3454
rect 132500 3460 132552 3466
rect 132500 3402 132552 3408
rect 134168 480 134196 4082
rect 135272 3534 135300 80022
rect 136652 4146 136680 80022
rect 136640 4140 136692 4146
rect 136640 4082 136692 4088
rect 138032 4078 138060 80022
rect 138020 4072 138072 4078
rect 138020 4014 138072 4020
rect 139412 4010 139440 80022
rect 140792 4826 140820 80022
rect 142172 6186 142200 80022
rect 142160 6180 142212 6186
rect 142160 6122 142212 6128
rect 140780 4820 140832 4826
rect 140780 4762 140832 4768
rect 139400 4004 139452 4010
rect 139400 3946 139452 3952
rect 143552 3942 143580 80022
rect 143540 3936 143592 3942
rect 143540 3878 143592 3884
rect 144932 3874 144960 80022
rect 144920 3868 144972 3874
rect 144920 3810 144972 3816
rect 146312 3806 146340 80022
rect 146300 3800 146352 3806
rect 146300 3742 146352 3748
rect 147692 3738 147720 80022
rect 147680 3732 147732 3738
rect 147680 3674 147732 3680
rect 149072 3670 149100 80022
rect 137652 3664 137704 3670
rect 137652 3606 137704 3612
rect 149060 3664 149112 3670
rect 149060 3606 149112 3612
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 137664 480 137692 3606
rect 150452 3602 150480 80022
rect 151832 16574 151860 80022
rect 151832 16546 151952 16574
rect 151820 4140 151872 4146
rect 151820 4082 151872 4088
rect 144736 3596 144788 3602
rect 144736 3538 144788 3544
rect 150440 3596 150492 3602
rect 150440 3538 150492 3544
rect 141240 3460 141292 3466
rect 141240 3402 141292 3408
rect 141252 480 141280 3402
rect 144748 480 144776 3538
rect 148324 3460 148376 3466
rect 148324 3402 148376 3408
rect 148336 480 148364 3402
rect 151832 480 151860 4082
rect 151924 3534 151952 16546
rect 151912 3528 151964 3534
rect 151912 3470 151964 3476
rect 153212 3466 153240 80022
rect 155420 77314 155448 80022
rect 156800 77314 156828 80022
rect 158180 77314 158208 80022
rect 159560 78198 159588 80022
rect 159548 78192 159600 78198
rect 159548 78134 159600 78140
rect 160940 78130 160968 80022
rect 160928 78124 160980 78130
rect 160928 78066 160980 78072
rect 162320 78062 162348 80022
rect 162308 78056 162360 78062
rect 162308 77998 162360 78004
rect 163700 77994 163728 80022
rect 163688 77988 163740 77994
rect 163688 77930 163740 77936
rect 155408 77308 155460 77314
rect 155408 77250 155460 77256
rect 156604 77308 156656 77314
rect 156604 77250 156656 77256
rect 156788 77308 156840 77314
rect 156788 77250 156840 77256
rect 157984 77308 158036 77314
rect 157984 77250 158036 77256
rect 158168 77308 158220 77314
rect 158168 77250 158220 77256
rect 159364 77308 159416 77314
rect 159364 77250 159416 77256
rect 156616 7614 156644 77250
rect 157996 10402 158024 77250
rect 159376 11762 159404 77250
rect 165080 75206 165108 80022
rect 165632 80022 166152 80050
rect 167012 80022 167532 80050
rect 168392 80022 168912 80050
rect 169772 80022 170292 80050
rect 171672 80022 172008 80050
rect 165068 75200 165120 75206
rect 165068 75142 165120 75148
rect 165632 13122 165660 80022
rect 167012 14482 167040 80022
rect 168392 43450 168420 80022
rect 168380 43444 168432 43450
rect 168380 43386 168432 43392
rect 169772 15910 169800 80022
rect 171980 77314 172008 80022
rect 172532 80022 173052 80050
rect 173912 80022 174432 80050
rect 175292 80022 175812 80050
rect 176672 80022 177192 80050
rect 178052 80022 178572 80050
rect 179432 80022 179952 80050
rect 180812 80022 181332 80050
rect 182192 80022 182712 80050
rect 183572 80022 184092 80050
rect 184952 80022 185472 80050
rect 186332 80022 186852 80050
rect 188232 80022 188568 80050
rect 189612 80022 189948 80050
rect 190992 80022 191328 80050
rect 192372 80022 192708 80050
rect 193752 80022 194088 80050
rect 195132 80022 195468 80050
rect 171968 77308 172020 77314
rect 171968 77250 172020 77256
rect 172532 18630 172560 80022
rect 173164 77308 173216 77314
rect 173164 77250 173216 77256
rect 172520 18624 172572 18630
rect 172520 18566 172572 18572
rect 169760 15904 169812 15910
rect 169760 15846 169812 15852
rect 167000 14476 167052 14482
rect 167000 14418 167052 14424
rect 165620 13116 165672 13122
rect 165620 13058 165672 13064
rect 159364 11756 159416 11762
rect 159364 11698 159416 11704
rect 157984 10396 158036 10402
rect 157984 10338 158036 10344
rect 173176 10334 173204 77250
rect 173164 10328 173216 10334
rect 173164 10270 173216 10276
rect 156604 7608 156656 7614
rect 156604 7550 156656 7556
rect 166080 6180 166132 6186
rect 166080 6122 166132 6128
rect 162492 4820 162544 4826
rect 162492 4762 162544 4768
rect 155408 4072 155460 4078
rect 155408 4014 155460 4020
rect 153200 3460 153252 3466
rect 153200 3402 153252 3408
rect 155420 480 155448 4014
rect 158904 4004 158956 4010
rect 158904 3946 158956 3952
rect 158916 480 158944 3946
rect 162504 480 162532 4762
rect 166092 480 166120 6122
rect 173912 5438 173940 80022
rect 173900 5432 173952 5438
rect 173900 5374 173952 5380
rect 175292 5370 175320 80022
rect 175280 5364 175332 5370
rect 175280 5306 175332 5312
rect 176672 5302 176700 80022
rect 176660 5296 176712 5302
rect 176660 5238 176712 5244
rect 178052 5234 178080 80022
rect 178040 5228 178092 5234
rect 178040 5170 178092 5176
rect 179432 5166 179460 80022
rect 179420 5160 179472 5166
rect 179420 5102 179472 5108
rect 180812 5098 180840 80022
rect 180800 5092 180852 5098
rect 180800 5034 180852 5040
rect 182192 5030 182220 80022
rect 182180 5024 182232 5030
rect 182180 4966 182232 4972
rect 183572 4962 183600 80022
rect 183560 4956 183612 4962
rect 183560 4898 183612 4904
rect 184952 4894 184980 80022
rect 184940 4888 184992 4894
rect 184940 4830 184992 4836
rect 186332 4826 186360 80022
rect 188540 78606 188568 80022
rect 188528 78600 188580 78606
rect 188528 78542 188580 78548
rect 189920 78538 189948 80022
rect 189908 78532 189960 78538
rect 189908 78474 189960 78480
rect 191300 78470 191328 80022
rect 191288 78464 191340 78470
rect 191288 78406 191340 78412
rect 192680 78402 192708 80022
rect 192668 78396 192720 78402
rect 192668 78338 192720 78344
rect 194060 78266 194088 80022
rect 195440 78334 195468 80022
rect 195992 80022 196512 80050
rect 197372 80022 197892 80050
rect 198752 80022 199272 80050
rect 200132 80022 200652 80050
rect 201512 80022 202032 80050
rect 202892 80022 203412 80050
rect 204272 80022 204792 80050
rect 205652 80022 206172 80050
rect 207032 80022 207552 80050
rect 208504 80022 208932 80050
rect 209792 80022 210312 80050
rect 211264 80022 211692 80050
rect 212552 80022 213072 80050
rect 214452 80022 214788 80050
rect 195428 78328 195480 78334
rect 195428 78270 195480 78276
rect 194048 78260 194100 78266
rect 194048 78202 194100 78208
rect 195992 73846 196020 80022
rect 195980 73840 196032 73846
rect 195980 73782 196032 73788
rect 197372 11830 197400 80022
rect 197360 11824 197412 11830
rect 197360 11766 197412 11772
rect 197912 7608 197964 7614
rect 197912 7550 197964 7556
rect 186320 4820 186372 4826
rect 186320 4762 186372 4768
rect 169576 3936 169628 3942
rect 169576 3878 169628 3884
rect 169588 480 169616 3878
rect 173164 3868 173216 3874
rect 173164 3810 173216 3816
rect 173176 480 173204 3810
rect 176660 3800 176712 3806
rect 176660 3742 176712 3748
rect 176672 480 176700 3742
rect 180248 3732 180300 3738
rect 180248 3674 180300 3680
rect 180260 480 180288 3674
rect 183744 3664 183796 3670
rect 183744 3606 183796 3612
rect 183756 480 183784 3606
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 187344 480 187372 3538
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 190840 480 190868 3470
rect 194416 3460 194468 3466
rect 194416 3402 194468 3408
rect 194428 480 194456 3402
rect 197924 480 197952 7550
rect 198752 6798 198780 80022
rect 199384 78600 199436 78606
rect 199384 78542 199436 78548
rect 198740 6792 198792 6798
rect 198740 6734 198792 6740
rect 199396 3534 199424 78542
rect 200132 6730 200160 80022
rect 200120 6724 200172 6730
rect 200120 6666 200172 6672
rect 201512 6662 201540 80022
rect 201592 10396 201644 10402
rect 201592 10338 201644 10344
rect 201500 6656 201552 6662
rect 201500 6598 201552 6604
rect 199384 3528 199436 3534
rect 201604 3482 201632 10338
rect 202892 6594 202920 80022
rect 203524 78532 203576 78538
rect 203524 78474 203576 78480
rect 202880 6588 202932 6594
rect 202880 6530 202932 6536
rect 203536 3806 203564 78474
rect 204272 6526 204300 80022
rect 205088 11756 205140 11762
rect 205088 11698 205140 11704
rect 204260 6520 204312 6526
rect 204260 6462 204312 6468
rect 203524 3800 203576 3806
rect 203524 3742 203576 3748
rect 199384 3470 199436 3476
rect 201512 3454 201632 3482
rect 201512 480 201540 3454
rect 205100 480 205128 11698
rect 205652 6458 205680 80022
rect 206284 78464 206336 78470
rect 206284 78406 206336 78412
rect 205640 6452 205692 6458
rect 205640 6394 205692 6400
rect 206296 3602 206324 78406
rect 207032 6390 207060 80022
rect 208400 78192 208452 78198
rect 208400 78134 208452 78140
rect 207020 6384 207072 6390
rect 207020 6326 207072 6332
rect 206284 3596 206336 3602
rect 206284 3538 206336 3544
rect 208412 3482 208440 78134
rect 208504 6322 208532 80022
rect 208492 6316 208544 6322
rect 208492 6258 208544 6264
rect 209792 6254 209820 80022
rect 210424 78396 210476 78402
rect 210424 78338 210476 78344
rect 209780 6248 209832 6254
rect 209780 6190 209832 6196
rect 210436 3738 210464 78338
rect 211160 78124 211212 78130
rect 211160 78066 211212 78072
rect 210424 3732 210476 3738
rect 210424 3674 210476 3680
rect 208412 3454 208624 3482
rect 208596 480 208624 3454
rect 211172 490 211200 78066
rect 211264 6186 211292 80022
rect 212552 44946 212580 80022
rect 214564 78328 214616 78334
rect 214564 78270 214616 78276
rect 213184 78260 213236 78266
rect 213184 78202 213236 78208
rect 212540 44940 212592 44946
rect 212540 44882 212592 44888
rect 211252 6180 211304 6186
rect 211252 6122 211304 6128
rect 213196 3670 213224 78202
rect 213184 3664 213236 3670
rect 213184 3606 213236 3612
rect 214576 3398 214604 78270
rect 214760 77314 214788 80022
rect 215404 80022 215832 80050
rect 216692 80022 217212 80050
rect 218592 80022 218928 80050
rect 215300 78056 215352 78062
rect 215300 77998 215352 78004
rect 214748 77308 214800 77314
rect 214748 77250 214800 77256
rect 214564 3392 214616 3398
rect 214564 3334 214616 3340
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211172 462 211752 490
rect 211724 354 211752 462
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 77998
rect 215404 36582 215432 80022
rect 215392 36576 215444 36582
rect 215392 36518 215444 36524
rect 216692 35222 216720 80022
rect 218900 77994 218928 80022
rect 219452 80022 219972 80050
rect 221352 80022 221688 80050
rect 218060 77988 218112 77994
rect 218060 77930 218112 77936
rect 218888 77988 218940 77994
rect 218888 77930 218940 77936
rect 217324 77308 217376 77314
rect 217324 77250 217376 77256
rect 216680 35216 216732 35222
rect 216680 35158 216732 35164
rect 217336 19990 217364 77250
rect 217324 19984 217376 19990
rect 217324 19926 217376 19932
rect 218072 3466 218100 77930
rect 219452 21486 219480 80022
rect 221660 77314 221688 80022
rect 222304 80022 222732 80050
rect 223592 80022 224112 80050
rect 225492 80022 225828 80050
rect 221648 77308 221700 77314
rect 221648 77250 221700 77256
rect 222200 75200 222252 75206
rect 222200 75142 222252 75148
rect 219440 21480 219492 21486
rect 219440 21422 219492 21428
rect 222212 16574 222240 75142
rect 222304 38010 222332 80022
rect 222292 38004 222344 38010
rect 222292 37946 222344 37952
rect 223592 25634 223620 80022
rect 225800 78674 225828 80022
rect 226352 80022 226872 80050
rect 227732 80022 228252 80050
rect 229112 80022 229632 80050
rect 230492 80022 231012 80050
rect 231872 80022 232392 80050
rect 233772 80022 234108 80050
rect 225788 78668 225840 78674
rect 225788 78610 225840 78616
rect 224224 77308 224276 77314
rect 224224 77250 224276 77256
rect 224236 49026 224264 77250
rect 224224 49020 224276 49026
rect 224224 48962 224276 48968
rect 226352 29714 226380 80022
rect 227732 43518 227760 80022
rect 228364 77988 228416 77994
rect 228364 77930 228416 77936
rect 227720 43512 227772 43518
rect 227720 43454 227772 43460
rect 226340 29708 226392 29714
rect 226340 29650 226392 29656
rect 223580 25628 223632 25634
rect 223580 25570 223632 25576
rect 228376 18698 228404 77930
rect 229112 31074 229140 80022
rect 230492 33794 230520 80022
rect 231124 78668 231176 78674
rect 231124 78610 231176 78616
rect 230480 33788 230532 33794
rect 230480 33730 230532 33736
rect 229100 31068 229152 31074
rect 229100 31010 229152 31016
rect 231136 26994 231164 78610
rect 231872 39438 231900 80022
rect 234080 78674 234108 80022
rect 234632 80022 235152 80050
rect 236532 80022 236868 80050
rect 234068 78668 234120 78674
rect 234068 78610 234120 78616
rect 233240 43444 233292 43450
rect 233240 43386 233292 43392
rect 231860 39432 231912 39438
rect 231860 39374 231912 39380
rect 231124 26988 231176 26994
rect 231124 26930 231176 26936
rect 228364 18692 228416 18698
rect 228364 18634 228416 18640
rect 233252 16574 233280 43386
rect 222212 16546 222792 16574
rect 233252 16546 233464 16574
rect 218060 3460 218112 3466
rect 218060 3402 218112 3408
rect 219256 3460 219308 3466
rect 219256 3402 219308 3408
rect 219268 480 219296 3402
rect 222764 480 222792 16546
rect 229376 14476 229428 14482
rect 229376 14418 229428 14424
rect 226340 13116 226392 13122
rect 226340 13058 226392 13064
rect 226352 480 226380 13058
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 14418
rect 233436 480 233464 16546
rect 234632 8158 234660 80022
rect 236840 78062 236868 80022
rect 237392 80022 237912 80050
rect 239292 80022 239628 80050
rect 240672 80022 241008 80050
rect 242052 80022 242388 80050
rect 236828 78056 236880 78062
rect 236828 77998 236880 78004
rect 236552 15904 236604 15910
rect 236552 15846 236604 15852
rect 234620 8152 234672 8158
rect 234620 8094 234672 8100
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 15846
rect 237392 8090 237420 80022
rect 239404 78668 239456 78674
rect 239404 78610 239456 78616
rect 239416 22846 239444 78610
rect 239600 77450 239628 80022
rect 239588 77444 239640 77450
rect 239588 77386 239640 77392
rect 240980 77314 241008 80022
rect 242164 78056 242216 78062
rect 242164 77998 242216 78004
rect 240968 77308 241020 77314
rect 240968 77250 241020 77256
rect 242176 24206 242204 77998
rect 242360 77382 242388 80022
rect 242912 80022 243432 80050
rect 244812 80022 245148 80050
rect 242348 77376 242400 77382
rect 242348 77318 242400 77324
rect 242256 77308 242308 77314
rect 242256 77250 242308 77256
rect 242268 44878 242296 77250
rect 242256 44872 242308 44878
rect 242256 44814 242308 44820
rect 242164 24200 242216 24206
rect 242164 24142 242216 24148
rect 239404 22840 239456 22846
rect 239404 22782 239456 22788
rect 240140 10328 240192 10334
rect 240140 10270 240192 10276
rect 237380 8084 237432 8090
rect 237380 8026 237432 8032
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 10270
rect 242912 8022 242940 80022
rect 244924 77444 244976 77450
rect 244924 77386 244976 77392
rect 244936 28354 244964 77386
rect 245120 77314 245148 80022
rect 245672 80022 246192 80050
rect 247572 80022 247908 80050
rect 245108 77308 245160 77314
rect 245108 77250 245160 77256
rect 245672 37942 245700 80022
rect 247880 77994 247908 80022
rect 248432 80022 248952 80050
rect 249812 80022 250332 80050
rect 251192 80022 251712 80050
rect 252572 80022 253092 80050
rect 253952 80022 254472 80050
rect 255852 80022 256188 80050
rect 247868 77988 247920 77994
rect 247868 77930 247920 77936
rect 246304 77376 246356 77382
rect 246304 77318 246356 77324
rect 245660 37936 245712 37942
rect 245660 37878 245712 37884
rect 244924 28348 244976 28354
rect 244924 28290 244976 28296
rect 242992 18624 243044 18630
rect 242992 18566 243044 18572
rect 243004 16574 243032 18566
rect 243004 16546 244136 16574
rect 242900 8016 242952 8022
rect 242900 7958 242952 7964
rect 244108 480 244136 16546
rect 246316 14550 246344 77318
rect 247684 77308 247736 77314
rect 247684 77250 247736 77256
rect 247696 17338 247724 77250
rect 247684 17332 247736 17338
rect 247684 17274 247736 17280
rect 246304 14544 246356 14550
rect 246304 14486 246356 14492
rect 248432 7954 248460 80022
rect 249812 13190 249840 80022
rect 249800 13184 249852 13190
rect 249800 13126 249852 13132
rect 248420 7948 248472 7954
rect 248420 7890 248472 7896
rect 251192 7886 251220 80022
rect 252572 10402 252600 80022
rect 252560 10396 252612 10402
rect 252560 10338 252612 10344
rect 251180 7880 251232 7886
rect 251180 7822 251232 7828
rect 253952 7818 253980 80022
rect 256160 78062 256188 80022
rect 256712 80022 257232 80050
rect 258092 80022 258612 80050
rect 259472 80022 259992 80050
rect 261372 80022 261708 80050
rect 256148 78056 256200 78062
rect 256148 77998 256200 78004
rect 253940 7812 253992 7818
rect 253940 7754 253992 7760
rect 256712 7750 256740 80022
rect 258092 15978 258120 80022
rect 258080 15972 258132 15978
rect 258080 15914 258132 15920
rect 256700 7744 256752 7750
rect 256700 7686 256752 7692
rect 259472 7682 259500 80022
rect 261680 78130 261708 80022
rect 262232 80022 262752 80050
rect 263612 80022 264132 80050
rect 264992 80022 265512 80050
rect 266372 80022 266892 80050
rect 267752 80022 268272 80050
rect 269132 80022 269652 80050
rect 270512 80022 271032 80050
rect 271892 80022 272412 80050
rect 273272 80022 273792 80050
rect 274652 80022 275172 80050
rect 276032 80022 276552 80050
rect 277412 80022 277932 80050
rect 278792 80022 279312 80050
rect 280172 80022 280692 80050
rect 281552 80022 282072 80050
rect 282932 80022 283452 80050
rect 284312 80022 284832 80050
rect 285692 80022 286212 80050
rect 287072 80022 287592 80050
rect 288452 80022 288972 80050
rect 289832 80022 290352 80050
rect 291212 80022 291732 80050
rect 292592 80022 293112 80050
rect 293972 80022 294492 80050
rect 295352 80022 295872 80050
rect 296732 80022 297252 80050
rect 298112 80022 298632 80050
rect 299492 80022 300012 80050
rect 300872 80022 301392 80050
rect 302252 80022 302772 80050
rect 304152 80022 304488 80050
rect 305532 80022 305868 80050
rect 306912 80022 307248 80050
rect 261668 78124 261720 78130
rect 261668 78066 261720 78072
rect 259460 7676 259512 7682
rect 259460 7618 259512 7624
rect 262232 7614 262260 80022
rect 263612 8974 263640 80022
rect 264992 40730 265020 80022
rect 264980 40724 265032 40730
rect 264980 40666 265032 40672
rect 266372 10334 266400 80022
rect 267752 11762 267780 80022
rect 269132 13122 269160 80022
rect 270512 14482 270540 80022
rect 271892 42090 271920 80022
rect 271880 42084 271932 42090
rect 271880 42026 271932 42032
rect 273272 15910 273300 80022
rect 274652 17270 274680 80022
rect 276032 28286 276060 80022
rect 276020 28280 276072 28286
rect 276020 28222 276072 28228
rect 274640 17264 274692 17270
rect 274640 17206 274692 17212
rect 273260 15904 273312 15910
rect 273260 15846 273312 15852
rect 270500 14476 270552 14482
rect 270500 14418 270552 14424
rect 269120 13116 269172 13122
rect 269120 13058 269172 13064
rect 267740 11756 267792 11762
rect 267740 11698 267792 11704
rect 266360 10328 266412 10334
rect 266360 10270 266412 10276
rect 263600 8968 263652 8974
rect 263600 8910 263652 8916
rect 262220 7608 262272 7614
rect 262220 7550 262272 7556
rect 277412 5438 277440 80022
rect 247592 5432 247644 5438
rect 247592 5374 247644 5380
rect 277400 5432 277452 5438
rect 277400 5374 277452 5380
rect 247604 480 247632 5374
rect 278792 5370 278820 80022
rect 251180 5364 251232 5370
rect 251180 5306 251232 5312
rect 278780 5364 278832 5370
rect 278780 5306 278832 5312
rect 251192 480 251220 5306
rect 280172 5302 280200 80022
rect 254676 5296 254728 5302
rect 254676 5238 254728 5244
rect 280160 5296 280212 5302
rect 280160 5238 280212 5244
rect 254688 480 254716 5238
rect 281552 5234 281580 80022
rect 258264 5228 258316 5234
rect 258264 5170 258316 5176
rect 281540 5228 281592 5234
rect 281540 5170 281592 5176
rect 258276 480 258304 5170
rect 282932 5166 282960 80022
rect 261760 5160 261812 5166
rect 261760 5102 261812 5108
rect 282920 5160 282972 5166
rect 282920 5102 282972 5108
rect 261772 480 261800 5102
rect 284312 5098 284340 80022
rect 265348 5092 265400 5098
rect 265348 5034 265400 5040
rect 284300 5092 284352 5098
rect 284300 5034 284352 5040
rect 265360 480 265388 5034
rect 285692 5030 285720 80022
rect 268844 5024 268896 5030
rect 268844 4966 268896 4972
rect 285680 5024 285732 5030
rect 285680 4966 285732 4972
rect 268856 480 268884 4966
rect 287072 4962 287100 80022
rect 272432 4956 272484 4962
rect 272432 4898 272484 4904
rect 287060 4956 287112 4962
rect 287060 4898 287112 4904
rect 272444 480 272472 4898
rect 288452 4894 288480 80022
rect 276020 4888 276072 4894
rect 276020 4830 276072 4836
rect 288440 4888 288492 4894
rect 288440 4830 288492 4836
rect 276032 480 276060 4830
rect 289832 4826 289860 80022
rect 291212 18630 291240 80022
rect 292592 24138 292620 80022
rect 292580 24132 292632 24138
rect 292580 24074 292632 24080
rect 293972 21418 294000 80022
rect 295352 22778 295380 80022
rect 296732 39370 296760 80022
rect 296720 39364 296772 39370
rect 296720 39306 296772 39312
rect 298112 25566 298140 80022
rect 299492 26926 299520 80022
rect 300872 43450 300900 80022
rect 300860 43444 300912 43450
rect 300860 43386 300912 43392
rect 302252 29646 302280 80022
rect 304460 78334 304488 80022
rect 304448 78328 304500 78334
rect 304448 78270 304500 78276
rect 305840 78198 305868 80022
rect 307220 78266 307248 80022
rect 307772 80022 308292 80050
rect 309152 80022 309672 80050
rect 311052 80022 311388 80050
rect 312432 80022 312768 80050
rect 315192 80022 315528 80050
rect 317952 80022 318288 80050
rect 307208 78260 307260 78266
rect 307208 78202 307260 78208
rect 305828 78192 305880 78198
rect 305828 78134 305880 78140
rect 303620 73840 303672 73846
rect 303620 73782 303672 73788
rect 302240 29640 302292 29646
rect 302240 29582 302292 29588
rect 299480 26920 299532 26926
rect 299480 26862 299532 26868
rect 298100 25560 298152 25566
rect 298100 25502 298152 25508
rect 295340 22772 295392 22778
rect 295340 22714 295392 22720
rect 293960 21412 294012 21418
rect 293960 21354 294012 21360
rect 291200 18624 291252 18630
rect 291200 18566 291252 18572
rect 303632 16574 303660 73782
rect 307772 48210 307800 80022
rect 309152 48278 309180 80022
rect 311360 78470 311388 80022
rect 312740 78674 312768 80022
rect 312728 78668 312780 78674
rect 312728 78610 312780 78616
rect 315500 78538 315528 80022
rect 318260 78742 318288 80022
rect 318248 78736 318300 78742
rect 318248 78678 318300 78684
rect 318352 78674 318380 93826
rect 318340 78668 318392 78674
rect 318340 78610 318392 78616
rect 319456 78538 319484 231814
rect 319536 230512 319588 230518
rect 319536 230454 319588 230460
rect 315488 78532 315540 78538
rect 315488 78474 315540 78480
rect 319444 78532 319496 78538
rect 319444 78474 319496 78480
rect 319548 78470 319576 230454
rect 358832 78742 358860 439175
rect 358924 353938 358952 596226
rect 359016 357882 359044 596838
rect 359096 596760 359148 596766
rect 359096 596702 359148 596708
rect 359108 358601 359136 596702
rect 359188 596556 359240 596562
rect 359188 596498 359240 596504
rect 359094 358592 359150 358601
rect 359094 358527 359150 358536
rect 359200 358426 359228 596498
rect 359738 560280 359794 560289
rect 359738 560215 359794 560224
rect 359752 559201 359780 560215
rect 359738 559192 359794 559201
rect 359738 559127 359794 559136
rect 359648 476944 359700 476950
rect 359648 476886 359700 476892
rect 359372 476808 359424 476814
rect 359372 476750 359424 476756
rect 359280 476196 359332 476202
rect 359280 476138 359332 476144
rect 359188 358420 359240 358426
rect 359188 358362 359240 358368
rect 359004 357876 359056 357882
rect 359004 357818 359056 357824
rect 359292 355366 359320 476138
rect 359384 358018 359412 476750
rect 359556 476740 359608 476746
rect 359556 476682 359608 476688
rect 359464 476604 359516 476610
rect 359464 476546 359516 476552
rect 359476 358358 359504 476546
rect 359568 358562 359596 476682
rect 359660 359446 359688 476886
rect 359752 454782 359780 559127
rect 360200 476400 360252 476406
rect 360200 476342 360252 476348
rect 359740 454776 359792 454782
rect 359740 454718 359792 454724
rect 359648 359440 359700 359446
rect 359648 359382 359700 359388
rect 359556 358556 359608 358562
rect 359556 358498 359608 358504
rect 359464 358352 359516 358358
rect 359464 358294 359516 358300
rect 359372 358012 359424 358018
rect 359372 357954 359424 357960
rect 360212 355570 360240 476342
rect 360292 476332 360344 476338
rect 360292 476274 360344 476280
rect 360200 355564 360252 355570
rect 360200 355506 360252 355512
rect 360304 355502 360332 476274
rect 360292 355496 360344 355502
rect 360292 355438 360344 355444
rect 359280 355360 359332 355366
rect 359280 355302 359332 355308
rect 358912 353932 358964 353938
rect 358912 353874 358964 353880
rect 360856 333266 360884 700334
rect 363604 700324 363656 700330
rect 363604 700266 363656 700272
rect 361672 476264 361724 476270
rect 361672 476206 361724 476212
rect 361580 359848 361632 359854
rect 361580 359790 361632 359796
rect 360844 333260 360896 333266
rect 360844 333202 360896 333208
rect 358820 78736 358872 78742
rect 358820 78678 358872 78684
rect 311348 78464 311400 78470
rect 311348 78406 311400 78412
rect 319536 78464 319588 78470
rect 319536 78406 319588 78412
rect 327724 78328 327776 78334
rect 327724 78270 327776 78276
rect 323584 78124 323636 78130
rect 323584 78066 323636 78072
rect 320824 78056 320876 78062
rect 320824 77998 320876 78004
rect 313924 77988 313976 77994
rect 313924 77930 313976 77936
rect 309140 48272 309192 48278
rect 309140 48214 309192 48220
rect 307760 48204 307812 48210
rect 307760 48146 307812 48152
rect 303632 16546 303936 16574
rect 279516 4820 279568 4826
rect 279516 4762 279568 4768
rect 289820 4820 289872 4826
rect 289820 4762 289872 4768
rect 279528 480 279556 4762
rect 286600 3800 286652 3806
rect 286600 3742 286652 3748
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 283116 480 283144 3470
rect 286612 480 286640 3742
rect 293684 3732 293736 3738
rect 293684 3674 293736 3680
rect 290188 3596 290240 3602
rect 290188 3538 290240 3544
rect 290200 480 290228 3538
rect 293696 480 293724 3674
rect 297272 3664 297324 3670
rect 297272 3606 297324 3612
rect 297284 480 297312 3606
rect 300768 3460 300820 3466
rect 300768 3402 300820 3408
rect 300780 480 300808 3402
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 307944 11824 307996 11830
rect 307944 11766 307996 11772
rect 307956 480 307984 11766
rect 311440 6792 311492 6798
rect 311440 6734 311492 6740
rect 311452 480 311480 6734
rect 313936 3806 313964 77930
rect 315028 6724 315080 6730
rect 315028 6666 315080 6672
rect 313924 3800 313976 3806
rect 313924 3742 313976 3748
rect 315040 480 315068 6666
rect 318524 6656 318576 6662
rect 318524 6598 318576 6604
rect 318536 480 318564 6598
rect 320836 3738 320864 77998
rect 322112 6588 322164 6594
rect 322112 6530 322164 6536
rect 320824 3732 320876 3738
rect 320824 3674 320876 3680
rect 322124 480 322152 6530
rect 323596 3670 323624 78066
rect 325608 6520 325660 6526
rect 325608 6462 325660 6468
rect 323584 3664 323636 3670
rect 323584 3606 323636 3612
rect 325620 480 325648 6462
rect 327736 3466 327764 78270
rect 331864 78260 331916 78266
rect 331864 78202 331916 78208
rect 330484 78192 330536 78198
rect 330484 78134 330536 78140
rect 329196 6452 329248 6458
rect 329196 6394 329248 6400
rect 327724 3460 327776 3466
rect 327724 3402 327776 3408
rect 329208 480 329236 6394
rect 330496 3602 330524 78134
rect 330484 3596 330536 3602
rect 330484 3538 330536 3544
rect 331876 3534 331904 78202
rect 361592 48210 361620 359790
rect 361684 355434 361712 476206
rect 362224 367192 362276 367198
rect 362224 367134 362276 367140
rect 362236 359854 362264 367134
rect 362224 359848 362276 359854
rect 362224 359790 362276 359796
rect 361672 355428 361724 355434
rect 361672 355370 361724 355376
rect 363616 319462 363644 700266
rect 364352 330546 364380 702406
rect 392584 700528 392636 700534
rect 392584 700470 392636 700476
rect 366364 700460 366416 700466
rect 366364 700402 366416 700408
rect 364340 330540 364392 330546
rect 364340 330482 364392 330488
rect 366376 324970 366404 700402
rect 378784 685908 378836 685914
rect 378784 685850 378836 685856
rect 378796 607918 378824 685850
rect 378784 607912 378836 607918
rect 378784 607854 378836 607860
rect 389822 597272 389878 597281
rect 389822 597207 389878 597216
rect 387524 594652 387576 594658
rect 387524 594594 387576 594600
rect 387156 594584 387208 594590
rect 387156 594526 387208 594532
rect 387064 594244 387116 594250
rect 387064 594186 387116 594192
rect 386972 594108 387024 594114
rect 386972 594050 387024 594056
rect 384396 591456 384448 591462
rect 384396 591398 384448 591404
rect 384304 591388 384356 591394
rect 384304 591330 384356 591336
rect 374644 487824 374696 487830
rect 374644 487766 374696 487772
rect 370502 477184 370558 477193
rect 370502 477119 370558 477128
rect 366364 324964 366416 324970
rect 366364 324906 366416 324912
rect 363604 319456 363656 319462
rect 363604 319398 363656 319404
rect 370516 312594 370544 477119
rect 374656 447098 374684 487766
rect 374644 447092 374696 447098
rect 374644 447034 374696 447040
rect 384316 348566 384344 591330
rect 384304 348560 384356 348566
rect 384304 348502 384356 348508
rect 384408 348498 384436 591398
rect 384488 591320 384540 591326
rect 384488 591262 384540 591268
rect 384500 348634 384528 591262
rect 384488 348628 384540 348634
rect 384488 348570 384540 348576
rect 384396 348492 384448 348498
rect 384396 348434 384448 348440
rect 386984 348226 387012 594050
rect 387076 348362 387104 594186
rect 387168 348838 387196 594526
rect 387340 594516 387392 594522
rect 387340 594458 387392 594464
rect 387248 594312 387300 594318
rect 387248 594254 387300 594260
rect 387260 349110 387288 594254
rect 387248 349104 387300 349110
rect 387248 349046 387300 349052
rect 387352 348906 387380 594458
rect 387432 594380 387484 594386
rect 387432 594322 387484 594328
rect 387444 349042 387472 594322
rect 387432 349036 387484 349042
rect 387432 348978 387484 348984
rect 387340 348900 387392 348906
rect 387340 348842 387392 348848
rect 387156 348832 387208 348838
rect 387156 348774 387208 348780
rect 387536 348770 387564 594594
rect 387616 594448 387668 594454
rect 387616 594390 387668 594396
rect 387628 348974 387656 594390
rect 387708 594176 387760 594182
rect 387708 594118 387760 594124
rect 387616 348968 387668 348974
rect 387616 348910 387668 348916
rect 387524 348764 387576 348770
rect 387524 348706 387576 348712
rect 387064 348356 387116 348362
rect 387064 348298 387116 348304
rect 387720 348294 387748 594118
rect 389730 594008 389786 594017
rect 389730 593943 389786 593952
rect 389744 351762 389772 593943
rect 389732 351756 389784 351762
rect 389732 351698 389784 351704
rect 389836 351490 389864 597207
rect 390192 594788 390244 594794
rect 390192 594730 390244 594736
rect 389916 594720 389968 594726
rect 389916 594662 389968 594668
rect 389824 351484 389876 351490
rect 389824 351426 389876 351432
rect 389928 348702 389956 594662
rect 390098 594416 390154 594425
rect 390098 594351 390154 594360
rect 390008 593972 390060 593978
rect 390008 593914 390060 593920
rect 390020 351830 390048 593914
rect 390008 351824 390060 351830
rect 390008 351766 390060 351772
rect 390112 351558 390140 594351
rect 390100 351552 390152 351558
rect 390100 351494 390152 351500
rect 390204 351150 390232 594730
rect 390466 594280 390522 594289
rect 390466 594215 390522 594224
rect 390282 594144 390338 594153
rect 390282 594079 390338 594088
rect 390296 351694 390324 594079
rect 390376 594040 390428 594046
rect 390376 593982 390428 593988
rect 390388 351898 390416 593982
rect 390376 351892 390428 351898
rect 390376 351834 390428 351840
rect 390284 351688 390336 351694
rect 390284 351630 390336 351636
rect 390480 351626 390508 594215
rect 392400 474156 392452 474162
rect 392400 474098 392452 474104
rect 392412 354482 392440 474098
rect 392492 471504 392544 471510
rect 392492 471446 392544 471452
rect 392400 354476 392452 354482
rect 392400 354418 392452 354424
rect 390468 351620 390520 351626
rect 390468 351562 390520 351568
rect 392504 351218 392532 471446
rect 392492 351212 392544 351218
rect 392492 351154 392544 351160
rect 390192 351144 390244 351150
rect 390192 351086 390244 351092
rect 389916 348696 389968 348702
rect 389916 348638 389968 348644
rect 387708 348288 387760 348294
rect 387708 348230 387760 348236
rect 386972 348220 387024 348226
rect 386972 348162 387024 348168
rect 392596 341562 392624 700470
rect 397472 699825 397500 703520
rect 413664 700466 413692 703520
rect 429856 700534 429884 703520
rect 429844 700528 429896 700534
rect 429844 700470 429896 700476
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 462332 700398 462360 703520
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 478524 700330 478552 703520
rect 494808 700505 494836 703520
rect 494794 700496 494850 700505
rect 494794 700431 494850 700440
rect 527192 700369 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 527178 700360 527234 700369
rect 478512 700324 478564 700330
rect 527178 700295 527234 700304
rect 478512 700266 478564 700272
rect 397458 699816 397514 699825
rect 397458 699751 397514 699760
rect 530950 685944 531006 685953
rect 530950 685879 530952 685888
rect 531004 685879 531006 685888
rect 536840 685908 536892 685914
rect 530952 685850 531004 685856
rect 536840 685850 536892 685856
rect 397274 636848 397330 636857
rect 397274 636783 397330 636792
rect 396906 635896 396962 635905
rect 396906 635831 396962 635840
rect 396630 632768 396686 632777
rect 396630 632703 396686 632712
rect 394700 607912 394752 607918
rect 394700 607854 394752 607860
rect 394712 607238 394740 607854
rect 394700 607232 394752 607238
rect 394700 607174 394752 607180
rect 392674 597408 392730 597417
rect 392674 597343 392730 597352
rect 392688 351393 392716 597343
rect 392858 596456 392914 596465
rect 392858 596391 392914 596400
rect 392768 471368 392820 471374
rect 392768 471310 392820 471316
rect 392674 351384 392730 351393
rect 392780 351354 392808 471310
rect 392872 351422 392900 596391
rect 394712 567186 394740 607174
rect 395344 597304 395396 597310
rect 395344 597246 395396 597252
rect 395068 593904 395120 593910
rect 395068 593846 395120 593852
rect 394700 567180 394752 567186
rect 394700 567122 394752 567128
rect 394332 477964 394384 477970
rect 394332 477906 394384 477912
rect 394056 476264 394108 476270
rect 394056 476206 394108 476212
rect 393964 474700 394016 474706
rect 393964 474642 394016 474648
rect 393044 474088 393096 474094
rect 393044 474030 393096 474036
rect 392952 474020 393004 474026
rect 392952 473962 393004 473968
rect 392964 354618 392992 473962
rect 392952 354612 393004 354618
rect 392952 354554 393004 354560
rect 393056 354550 393084 474030
rect 393228 471436 393280 471442
rect 393228 471378 393280 471384
rect 393136 471300 393188 471306
rect 393136 471242 393188 471248
rect 393044 354544 393096 354550
rect 393044 354486 393096 354492
rect 392860 351416 392912 351422
rect 392860 351358 392912 351364
rect 392674 351319 392730 351328
rect 392768 351348 392820 351354
rect 392768 351290 392820 351296
rect 393148 351014 393176 471242
rect 393240 351286 393268 471378
rect 393872 471232 393924 471238
rect 393872 471174 393924 471180
rect 393780 359848 393832 359854
rect 393780 359790 393832 359796
rect 393792 356522 393820 359790
rect 393884 356561 393912 471174
rect 393976 356697 394004 474642
rect 394068 357134 394096 476206
rect 394148 476196 394200 476202
rect 394148 476138 394200 476144
rect 394160 359854 394188 476138
rect 394240 476128 394292 476134
rect 394240 476070 394292 476076
rect 394148 359848 394200 359854
rect 394148 359790 394200 359796
rect 394252 359530 394280 476070
rect 394160 359502 394280 359530
rect 394056 357128 394108 357134
rect 394056 357070 394108 357076
rect 393962 356688 394018 356697
rect 393962 356623 394018 356632
rect 394160 356590 394188 359502
rect 394344 359394 394372 477906
rect 394424 477896 394476 477902
rect 394424 477838 394476 477844
rect 394252 359366 394372 359394
rect 394252 357270 394280 359366
rect 394436 359258 394464 477838
rect 394516 477760 394568 477766
rect 394516 477702 394568 477708
rect 394344 359230 394464 359258
rect 394240 357264 394292 357270
rect 394240 357206 394292 357212
rect 394252 356590 394280 357206
rect 394344 356930 394372 359230
rect 394424 357128 394476 357134
rect 394424 357070 394476 357076
rect 394332 356924 394384 356930
rect 394332 356866 394384 356872
rect 394436 356658 394464 357070
rect 394528 356794 394556 477702
rect 394608 477692 394660 477698
rect 394608 477634 394660 477640
rect 394620 357066 394648 477634
rect 395080 474706 395108 593846
rect 395160 591524 395212 591530
rect 395160 591466 395212 591472
rect 395068 474700 395120 474706
rect 395068 474642 395120 474648
rect 395080 473822 395108 474642
rect 395068 473816 395120 473822
rect 395068 473758 395120 473764
rect 395172 471986 395200 591466
rect 395252 474292 395304 474298
rect 395252 474234 395304 474240
rect 395160 471980 395212 471986
rect 395160 471922 395212 471928
rect 395172 471238 395200 471922
rect 395160 471232 395212 471238
rect 395160 471174 395212 471180
rect 395264 359786 395292 474234
rect 395252 359780 395304 359786
rect 395252 359722 395304 359728
rect 394608 357060 394660 357066
rect 394608 357002 394660 357008
rect 394608 356924 394660 356930
rect 394608 356866 394660 356872
rect 394516 356788 394568 356794
rect 394516 356730 394568 356736
rect 394514 356688 394570 356697
rect 394424 356652 394476 356658
rect 394620 356658 394648 356866
rect 394514 356623 394570 356632
rect 394608 356652 394660 356658
rect 394424 356594 394476 356600
rect 394148 356584 394200 356590
rect 393870 356552 393926 356561
rect 393780 356516 393832 356522
rect 394148 356526 394200 356532
rect 394240 356584 394292 356590
rect 394240 356526 394292 356532
rect 393870 356487 393926 356496
rect 393780 356458 393832 356464
rect 394160 356182 394188 356526
rect 394528 356425 394556 356623
rect 394608 356594 394660 356600
rect 394608 356516 394660 356522
rect 394608 356458 394660 356464
rect 394514 356416 394570 356425
rect 394514 356351 394570 356360
rect 394148 356176 394200 356182
rect 394148 356118 394200 356124
rect 394620 356114 394648 356458
rect 394608 356108 394660 356114
rect 394608 356050 394660 356056
rect 393228 351280 393280 351286
rect 393228 351222 393280 351228
rect 393136 351008 393188 351014
rect 393136 350950 393188 350956
rect 392584 341556 392636 341562
rect 392584 341498 392636 341504
rect 395356 337482 395384 597246
rect 395804 591592 395856 591598
rect 395804 591534 395856 591540
rect 395816 476610 395844 591534
rect 396446 516216 396502 516225
rect 396446 516151 396502 516160
rect 395804 476604 395856 476610
rect 395804 476546 395856 476552
rect 395816 476202 395844 476546
rect 395804 476196 395856 476202
rect 395804 476138 395856 476144
rect 395436 474700 395488 474706
rect 395436 474642 395488 474648
rect 395448 354074 395476 474642
rect 395620 474632 395672 474638
rect 395620 474574 395672 474580
rect 395528 473952 395580 473958
rect 395528 473894 395580 473900
rect 395436 354068 395488 354074
rect 395436 354010 395488 354016
rect 395540 354006 395568 473894
rect 395632 354142 395660 474574
rect 395712 474564 395764 474570
rect 395712 474506 395764 474512
rect 395724 354210 395752 474506
rect 395804 474496 395856 474502
rect 395804 474438 395856 474444
rect 395816 354278 395844 474438
rect 395988 474428 396040 474434
rect 395988 474370 396040 474376
rect 395896 474360 395948 474366
rect 395896 474302 395948 474308
rect 395908 354414 395936 474302
rect 395896 354408 395948 354414
rect 395896 354350 395948 354356
rect 396000 354346 396028 474370
rect 396460 454714 396488 516151
rect 396538 514856 396594 514865
rect 396538 514791 396594 514800
rect 396448 454708 396500 454714
rect 396448 454650 396500 454656
rect 396552 450566 396580 514791
rect 396644 512825 396672 632703
rect 396814 628144 396870 628153
rect 396814 628079 396870 628088
rect 396722 610056 396778 610065
rect 396722 609991 396778 610000
rect 396630 512816 396686 512825
rect 396630 512751 396686 512760
rect 396736 489977 396764 609991
rect 396828 508201 396856 628079
rect 396920 515953 396948 635831
rect 396998 633720 397054 633729
rect 396998 633655 397054 633664
rect 396906 515944 396962 515953
rect 396906 515879 396962 515888
rect 396920 514865 396948 515879
rect 396906 514856 396962 514865
rect 396906 514791 396962 514800
rect 397012 513777 397040 633655
rect 397090 631000 397146 631009
rect 397090 630935 397146 630944
rect 396998 513768 397054 513777
rect 396998 513703 397054 513712
rect 396998 512816 397054 512825
rect 396998 512751 397054 512760
rect 396906 510504 396962 510513
rect 396906 510439 396962 510448
rect 396920 509969 396948 510439
rect 396906 509960 396962 509969
rect 396906 509895 396962 509904
rect 396814 508192 396870 508201
rect 396814 508127 396870 508136
rect 396722 489968 396778 489977
rect 396722 489903 396778 489912
rect 396632 454708 396684 454714
rect 396632 454650 396684 454656
rect 396540 450560 396592 450566
rect 396540 450502 396592 450508
rect 396552 396001 396580 450502
rect 396644 396953 396672 454650
rect 396630 396944 396686 396953
rect 396630 396879 396686 396888
rect 396538 395992 396594 396001
rect 396538 395927 396594 395936
rect 396630 394632 396686 394641
rect 396630 394567 396686 394576
rect 396644 393825 396672 394567
rect 396630 393816 396686 393825
rect 396630 393751 396686 393760
rect 396446 370016 396502 370025
rect 396446 369951 396502 369960
rect 396460 367062 396488 369951
rect 396538 368112 396594 368121
rect 396538 368047 396594 368056
rect 396552 367130 396580 368047
rect 396540 367124 396592 367130
rect 396540 367066 396592 367072
rect 396448 367056 396500 367062
rect 396448 366998 396500 367004
rect 396644 360058 396672 393751
rect 396736 370025 396764 489903
rect 396828 388249 396856 508127
rect 396920 390017 396948 509895
rect 397012 392873 397040 512751
rect 397104 511057 397132 630935
rect 397182 608288 397238 608297
rect 397182 608223 397238 608232
rect 397196 607238 397224 608223
rect 397184 607232 397236 607238
rect 397184 607174 397236 607180
rect 397090 511048 397146 511057
rect 397090 510983 397146 510992
rect 396998 392864 397054 392873
rect 396998 392799 397054 392808
rect 396906 390008 396962 390017
rect 396906 389943 396962 389952
rect 396814 388240 396870 388249
rect 396814 388175 396870 388184
rect 396722 370016 396778 370025
rect 396722 369951 396778 369960
rect 396722 368384 396778 368393
rect 396722 368319 396778 368328
rect 396736 367198 396764 368319
rect 396724 367192 396776 367198
rect 396724 367134 396776 367140
rect 396724 367056 396776 367062
rect 396724 366998 396776 367004
rect 396632 360052 396684 360058
rect 396632 359994 396684 360000
rect 395988 354340 396040 354346
rect 395988 354282 396040 354288
rect 395804 354272 395856 354278
rect 395804 354214 395856 354220
rect 395712 354204 395764 354210
rect 395712 354146 395764 354152
rect 395620 354136 395672 354142
rect 395620 354078 395672 354084
rect 395528 354000 395580 354006
rect 395528 353942 395580 353948
rect 395344 337476 395396 337482
rect 395344 337418 395396 337424
rect 370504 312588 370556 312594
rect 370504 312530 370556 312536
rect 396736 289814 396764 366998
rect 396828 358766 396856 388175
rect 396816 358760 396868 358766
rect 396816 358702 396868 358708
rect 396920 358630 396948 389943
rect 396908 358624 396960 358630
rect 396908 358566 396960 358572
rect 397012 358086 397040 392799
rect 397104 391105 397132 510983
rect 397196 488345 397224 607174
rect 397288 516905 397316 636783
rect 397366 629912 397422 629921
rect 397366 629847 397422 629856
rect 397274 516896 397330 516905
rect 397274 516831 397330 516840
rect 397288 516225 397316 516831
rect 397274 516216 397330 516225
rect 397274 516151 397330 516160
rect 397380 510513 397408 629847
rect 435914 599584 435970 599593
rect 435914 599519 435970 599528
rect 415398 597544 415454 597553
rect 397736 597508 397788 597514
rect 415398 597479 415454 597488
rect 416778 597544 416834 597553
rect 416778 597479 416834 597488
rect 418158 597544 418214 597553
rect 418158 597479 418214 597488
rect 419538 597544 419594 597553
rect 419538 597479 419594 597488
rect 420918 597544 420974 597553
rect 420918 597479 420974 597488
rect 423126 597544 423182 597553
rect 423126 597479 423182 597488
rect 424966 597544 425022 597553
rect 424966 597479 425022 597488
rect 425610 597544 425666 597553
rect 425610 597479 425666 597488
rect 426530 597544 426586 597553
rect 426530 597479 426586 597488
rect 427634 597544 427690 597553
rect 427634 597479 427690 597488
rect 428002 597544 428058 597553
rect 428002 597479 428058 597488
rect 429198 597544 429254 597553
rect 429198 597479 429254 597488
rect 430578 597544 430634 597553
rect 430578 597479 430634 597488
rect 433338 597544 433394 597553
rect 433338 597479 433394 597488
rect 434534 597544 434590 597553
rect 434718 597544 434774 597553
rect 434590 597502 434668 597530
rect 434534 597479 434590 597488
rect 397736 597450 397788 597456
rect 397366 510504 397422 510513
rect 397366 510439 397422 510448
rect 397182 488336 397238 488345
rect 397182 488271 397238 488280
rect 397196 487830 397224 488271
rect 397184 487824 397236 487830
rect 397184 487766 397236 487772
rect 397196 487393 397224 487766
rect 397182 487384 397238 487393
rect 397182 487319 397238 487328
rect 397276 477828 397328 477834
rect 397276 477770 397328 477776
rect 397184 477624 397236 477630
rect 397184 477566 397236 477572
rect 397196 476814 397224 477566
rect 397184 476808 397236 476814
rect 397184 476750 397236 476756
rect 397090 391096 397146 391105
rect 397090 391031 397146 391040
rect 397104 358698 397132 391031
rect 397092 358692 397144 358698
rect 397092 358634 397144 358640
rect 397000 358080 397052 358086
rect 397000 358022 397052 358028
rect 397196 356833 397224 476750
rect 397288 359258 397316 477770
rect 397368 477556 397420 477562
rect 397368 477498 397420 477504
rect 397380 359378 397408 477498
rect 397748 476406 397776 597450
rect 399484 597440 399536 597446
rect 399484 597382 399536 597388
rect 397828 597372 397880 597378
rect 397828 597314 397880 597320
rect 397840 476542 397868 597314
rect 398288 596896 398340 596902
rect 398288 596838 398340 596844
rect 398104 596760 398156 596766
rect 398104 596702 398156 596708
rect 398012 592000 398064 592006
rect 398012 591942 398064 591948
rect 397920 591864 397972 591870
rect 397920 591806 397972 591812
rect 397932 478310 397960 591806
rect 398024 478446 398052 591942
rect 398012 478440 398064 478446
rect 398012 478382 398064 478388
rect 397920 478304 397972 478310
rect 397920 478246 397972 478252
rect 397932 477698 397960 478246
rect 398024 477766 398052 478382
rect 398012 477760 398064 477766
rect 398012 477702 398064 477708
rect 397920 477692 397972 477698
rect 397920 477634 397972 477640
rect 398116 477630 398144 596702
rect 398196 591796 398248 591802
rect 398196 591738 398248 591744
rect 398208 478242 398236 591738
rect 398196 478236 398248 478242
rect 398196 478178 398248 478184
rect 398104 477624 398156 477630
rect 398104 477566 398156 477572
rect 398208 477562 398236 478178
rect 398300 477766 398328 596838
rect 398564 596828 398616 596834
rect 398564 596770 398616 596776
rect 398472 596624 398524 596630
rect 398472 596566 398524 596572
rect 398380 596556 398432 596562
rect 398380 596498 398432 596504
rect 398392 478582 398420 596498
rect 398380 478576 398432 478582
rect 398380 478518 398432 478524
rect 398392 477970 398420 478518
rect 398380 477964 398432 477970
rect 398380 477906 398432 477912
rect 398288 477760 398340 477766
rect 398288 477702 398340 477708
rect 398484 477698 398512 596566
rect 398576 480254 398604 596770
rect 399300 591932 399352 591938
rect 399300 591874 399352 591880
rect 399208 591728 399260 591734
rect 399208 591670 399260 591676
rect 398576 480226 398788 480254
rect 398760 477714 398788 480226
rect 399220 478174 399248 591670
rect 399312 478378 399340 591874
rect 399392 591660 399444 591666
rect 399392 591602 399444 591608
rect 399300 478372 399352 478378
rect 399300 478314 399352 478320
rect 399208 478168 399260 478174
rect 399208 478110 399260 478116
rect 398472 477692 398524 477698
rect 398760 477686 398880 477714
rect 398472 477634 398524 477640
rect 398196 477556 398248 477562
rect 398196 477498 398248 477504
rect 398484 477442 398512 477634
rect 398748 477556 398800 477562
rect 398748 477498 398800 477504
rect 398484 477414 398696 477442
rect 398562 477320 398618 477329
rect 398562 477255 398618 477264
rect 398102 476640 398158 476649
rect 398102 476575 398158 476584
rect 397828 476536 397880 476542
rect 397828 476478 397880 476484
rect 397736 476400 397788 476406
rect 397736 476342 397788 476348
rect 397748 476270 397776 476342
rect 397736 476264 397788 476270
rect 397736 476206 397788 476212
rect 397840 476134 397868 476478
rect 397828 476128 397880 476134
rect 397828 476070 397880 476076
rect 397826 474328 397882 474337
rect 397826 474263 397882 474272
rect 397840 359650 397868 474263
rect 398010 474056 398066 474065
rect 398010 473991 398066 474000
rect 397920 473884 397972 473890
rect 397920 473826 397972 473832
rect 397828 359644 397880 359650
rect 397828 359586 397880 359592
rect 397368 359372 397420 359378
rect 397368 359314 397420 359320
rect 397288 359230 397408 359258
rect 397276 359168 397328 359174
rect 397276 359110 397328 359116
rect 397288 356930 397316 359110
rect 397380 357202 397408 359230
rect 397368 357196 397420 357202
rect 397368 357138 397420 357144
rect 397276 356924 397328 356930
rect 397276 356866 397328 356872
rect 397182 356824 397238 356833
rect 397182 356759 397238 356768
rect 397288 356318 397316 356866
rect 397380 356454 397408 357138
rect 397368 356448 397420 356454
rect 397368 356390 397420 356396
rect 397276 356312 397328 356318
rect 397276 356254 397328 356260
rect 397932 354385 397960 473826
rect 398024 359718 398052 473991
rect 398012 359712 398064 359718
rect 398012 359654 398064 359660
rect 397918 354376 397974 354385
rect 397918 354311 397974 354320
rect 398116 354113 398144 476575
rect 398286 476368 398342 476377
rect 398286 476303 398342 476312
rect 398194 474464 398250 474473
rect 398194 474399 398250 474408
rect 398208 359582 398236 474399
rect 398196 359576 398248 359582
rect 398196 359518 398248 359524
rect 398196 357332 398248 357338
rect 398196 357274 398248 357280
rect 398208 356726 398236 357274
rect 398196 356720 398248 356726
rect 398196 356662 398248 356668
rect 398300 354249 398328 476303
rect 398470 474192 398526 474201
rect 398470 474127 398526 474136
rect 398380 357060 398432 357066
rect 398380 357002 398432 357008
rect 398392 356386 398420 357002
rect 398380 356380 398432 356386
rect 398380 356322 398432 356328
rect 398484 354521 398512 474127
rect 398576 359514 398604 477255
rect 398564 359508 398616 359514
rect 398564 359450 398616 359456
rect 398668 357338 398696 477414
rect 398656 357332 398708 357338
rect 398656 357274 398708 357280
rect 398760 357066 398788 477498
rect 398852 476950 398880 477686
rect 399024 477624 399076 477630
rect 399024 477566 399076 477572
rect 398840 476944 398892 476950
rect 398840 476886 398892 476892
rect 398932 476264 398984 476270
rect 398932 476206 398984 476212
rect 398944 357377 398972 476206
rect 398930 357368 398986 357377
rect 398840 357332 398892 357338
rect 398930 357303 398986 357312
rect 398840 357274 398892 357280
rect 398748 357060 398800 357066
rect 398748 357002 398800 357008
rect 398852 356862 398880 357274
rect 398840 356856 398892 356862
rect 398840 356798 398892 356804
rect 398944 356289 398972 357303
rect 399036 357202 399064 477566
rect 399220 477562 399248 478110
rect 399312 477834 399340 478314
rect 399300 477828 399352 477834
rect 399300 477770 399352 477776
rect 399404 477562 399432 591602
rect 399496 477630 399524 597382
rect 399668 597032 399720 597038
rect 399668 596974 399720 596980
rect 399576 596488 399628 596494
rect 399576 596430 399628 596436
rect 399588 478514 399616 596430
rect 399576 478508 399628 478514
rect 399576 478450 399628 478456
rect 399588 477902 399616 478450
rect 399576 477896 399628 477902
rect 399576 477838 399628 477844
rect 399484 477624 399536 477630
rect 399484 477566 399536 477572
rect 399208 477556 399260 477562
rect 399208 477498 399260 477504
rect 399392 477556 399444 477562
rect 399392 477498 399444 477504
rect 399404 476354 399432 477498
rect 399680 477222 399708 596974
rect 399944 596964 399996 596970
rect 399944 596906 399996 596912
rect 399760 596692 399812 596698
rect 399760 596634 399812 596640
rect 399668 477216 399720 477222
rect 399668 477158 399720 477164
rect 399484 477012 399536 477018
rect 399484 476954 399536 476960
rect 399128 476326 399432 476354
rect 399128 357338 399156 476326
rect 399208 476196 399260 476202
rect 399208 476138 399260 476144
rect 399220 358154 399248 476138
rect 399300 476128 399352 476134
rect 399300 476070 399352 476076
rect 399208 358148 399260 358154
rect 399208 358090 399260 358096
rect 399312 357406 399340 476070
rect 399496 475946 399524 476954
rect 399576 476944 399628 476950
rect 399576 476886 399628 476892
rect 399404 475918 399524 475946
rect 399300 357400 399352 357406
rect 399300 357342 399352 357348
rect 399116 357332 399168 357338
rect 399116 357274 399168 357280
rect 399404 357241 399432 475918
rect 399484 474224 399536 474230
rect 399484 474166 399536 474172
rect 399390 357232 399446 357241
rect 399024 357196 399076 357202
rect 399390 357167 399446 357176
rect 399024 357138 399076 357144
rect 398930 356280 398986 356289
rect 399036 356250 399064 357138
rect 398930 356215 398986 356224
rect 399024 356244 399076 356250
rect 399024 356186 399076 356192
rect 398470 354512 398526 354521
rect 398470 354447 398526 354456
rect 398286 354240 398342 354249
rect 398286 354175 398342 354184
rect 398102 354104 398158 354113
rect 398102 354039 398158 354048
rect 399496 351082 399524 474166
rect 399588 357105 399616 476886
rect 399680 476270 399708 477158
rect 399772 476882 399800 596634
rect 399852 596216 399904 596222
rect 399852 596158 399904 596164
rect 399864 477154 399892 596158
rect 399852 477148 399904 477154
rect 399852 477090 399904 477096
rect 399760 476876 399812 476882
rect 399760 476818 399812 476824
rect 399668 476264 399720 476270
rect 399668 476206 399720 476212
rect 399772 476134 399800 476818
rect 399864 476202 399892 477090
rect 399956 477086 399984 596906
rect 415412 596222 415440 597479
rect 416792 597038 416820 597479
rect 416780 597032 416832 597038
rect 416780 596974 416832 596980
rect 418172 596902 418200 597479
rect 419552 596970 419580 597479
rect 419540 596964 419592 596970
rect 419540 596906 419592 596912
rect 418160 596896 418212 596902
rect 418160 596838 418212 596844
rect 419540 596828 419592 596834
rect 419540 596770 419592 596776
rect 419552 596737 419580 596770
rect 420932 596766 420960 597479
rect 423140 596834 423168 597479
rect 424980 597106 425008 597479
rect 425624 597174 425652 597479
rect 426544 597242 426572 597479
rect 426532 597236 426584 597242
rect 426532 597178 426584 597184
rect 425612 597168 425664 597174
rect 425612 597110 425664 597116
rect 424968 597100 425020 597106
rect 424968 597042 425020 597048
rect 423128 596828 423180 596834
rect 423128 596770 423180 596776
rect 420920 596760 420972 596766
rect 419538 596728 419594 596737
rect 420920 596702 420972 596708
rect 419538 596663 419594 596672
rect 424980 596630 425008 597042
rect 424968 596624 425020 596630
rect 424968 596566 425020 596572
rect 425624 596562 425652 597110
rect 425612 596556 425664 596562
rect 425612 596498 425664 596504
rect 426440 596556 426492 596562
rect 426440 596498 426492 596504
rect 415400 596216 415452 596222
rect 415400 596158 415452 596164
rect 426452 592006 426480 596498
rect 426544 596494 426572 597178
rect 427648 596562 427676 597479
rect 427818 596728 427874 596737
rect 427818 596663 427874 596672
rect 427636 596556 427688 596562
rect 427636 596498 427688 596504
rect 426532 596488 426584 596494
rect 426532 596430 426584 596436
rect 426440 592000 426492 592006
rect 426440 591942 426492 591948
rect 427832 571985 427860 596663
rect 428016 596630 428044 597479
rect 428004 596624 428056 596630
rect 428004 596566 428056 596572
rect 428016 591870 428044 596566
rect 429212 596494 429240 597479
rect 429200 596488 429252 596494
rect 429200 596430 429252 596436
rect 429212 591938 429240 596430
rect 429200 591932 429252 591938
rect 429200 591874 429252 591880
rect 428004 591864 428056 591870
rect 428004 591806 428056 591812
rect 427818 571976 427874 571985
rect 427818 571911 427874 571920
rect 430592 570625 430620 597479
rect 430670 596728 430726 596737
rect 430670 596663 430726 596672
rect 431958 596728 432014 596737
rect 431958 596663 432014 596672
rect 430684 596290 430712 596663
rect 431972 596426 432000 596663
rect 431960 596420 432012 596426
rect 431960 596362 432012 596368
rect 430672 596284 430724 596290
rect 430672 596226 430724 596232
rect 430684 591802 430712 596226
rect 430672 591796 430724 591802
rect 430672 591738 430724 591744
rect 431972 591734 432000 596362
rect 431960 591728 432012 591734
rect 431960 591670 432012 591676
rect 430578 570616 430634 570625
rect 430578 570551 430634 570560
rect 433352 563689 433380 597479
rect 434640 597446 434668 597502
rect 435928 597530 435956 599519
rect 451094 599448 451150 599457
rect 451094 599383 451150 599392
rect 437110 597544 437166 597553
rect 435928 597514 436048 597530
rect 435928 597508 436060 597514
rect 435928 597502 436008 597508
rect 434718 597479 434774 597488
rect 434628 597440 434680 597446
rect 434628 597382 434680 597388
rect 434640 597038 434668 597382
rect 434732 597310 434760 597479
rect 437110 597479 437166 597488
rect 437478 597544 437534 597553
rect 437478 597479 437534 597488
rect 438858 597544 438914 597553
rect 438858 597479 438914 597488
rect 441986 597544 442042 597553
rect 441986 597479 442042 597488
rect 442998 597544 443054 597553
rect 442998 597479 443054 597488
rect 443642 597544 443698 597553
rect 443642 597479 443698 597488
rect 444378 597544 444434 597553
rect 444378 597479 444434 597488
rect 445758 597544 445814 597553
rect 445758 597479 445814 597488
rect 447138 597544 447194 597553
rect 447138 597479 447194 597488
rect 449898 597544 449954 597553
rect 449898 597479 449954 597488
rect 436008 597450 436060 597456
rect 434720 597304 434772 597310
rect 434720 597246 434772 597252
rect 434628 597032 434680 597038
rect 434628 596974 434680 596980
rect 436020 596970 436048 597450
rect 437124 597378 437152 597479
rect 437112 597372 437164 597378
rect 437112 597314 437164 597320
rect 436008 596964 436060 596970
rect 436008 596906 436060 596912
rect 437124 596902 437152 597314
rect 437112 596896 437164 596902
rect 437112 596838 437164 596844
rect 433430 596728 433486 596737
rect 433430 596663 433486 596672
rect 433444 596358 433472 596663
rect 433432 596352 433484 596358
rect 433432 596294 433484 596300
rect 433444 591666 433472 596294
rect 437492 596222 437520 597479
rect 438872 596737 438900 597479
rect 440330 597136 440386 597145
rect 442000 597106 442028 597479
rect 440330 597071 440386 597080
rect 441988 597100 442040 597106
rect 438858 596728 438914 596737
rect 438858 596663 438914 596672
rect 437480 596216 437532 596222
rect 437480 596158 437532 596164
rect 433432 591660 433484 591666
rect 433432 591602 433484 591608
rect 437492 591598 437520 596158
rect 438872 593910 438900 596663
rect 438860 593904 438912 593910
rect 438860 593846 438912 593852
rect 437480 591592 437532 591598
rect 437480 591534 437532 591540
rect 440344 591530 440372 597071
rect 441988 597042 442040 597048
rect 441618 597000 441674 597009
rect 441618 596935 441674 596944
rect 441632 596834 441660 596935
rect 441620 596828 441672 596834
rect 441620 596770 441672 596776
rect 443012 594561 443040 597479
rect 443656 597174 443684 597479
rect 444392 597242 444420 597479
rect 444380 597236 444432 597242
rect 444380 597178 444432 597184
rect 443644 597168 443696 597174
rect 443644 597110 443696 597116
rect 442998 594552 443054 594561
rect 442998 594487 443054 594496
rect 440332 591524 440384 591530
rect 440332 591466 440384 591472
rect 445772 591462 445800 597479
rect 445850 597000 445906 597009
rect 445850 596935 445906 596944
rect 445864 596562 445892 596935
rect 445852 596556 445904 596562
rect 445852 596498 445904 596504
rect 445760 591456 445812 591462
rect 445760 591398 445812 591404
rect 447152 591394 447180 597479
rect 447230 597000 447286 597009
rect 447230 596935 447286 596944
rect 448518 597000 448574 597009
rect 448518 596935 448574 596944
rect 447244 596630 447272 596935
rect 447232 596624 447284 596630
rect 447232 596566 447284 596572
rect 448532 596494 448560 596935
rect 448520 596488 448572 596494
rect 448520 596430 448572 596436
rect 448518 596320 448574 596329
rect 448518 596255 448520 596264
rect 448572 596255 448574 596264
rect 448520 596226 448572 596232
rect 447140 591388 447192 591394
rect 447140 591330 447192 591336
rect 449912 591326 449940 597479
rect 451108 596465 451136 599383
rect 462318 597544 462374 597553
rect 462318 597479 462374 597488
rect 465078 597544 465134 597553
rect 465078 597479 465134 597488
rect 467838 597544 467894 597553
rect 467838 597479 467894 597488
rect 473358 597544 473414 597553
rect 473358 597479 473414 597488
rect 474738 597544 474794 597553
rect 474738 597479 474794 597488
rect 477498 597544 477554 597553
rect 477498 597479 477554 597488
rect 483018 597544 483074 597553
rect 483018 597479 483074 597488
rect 485778 597544 485834 597553
rect 485778 597479 485834 597488
rect 488538 597544 488594 597553
rect 488538 597479 488594 597488
rect 495438 597544 495494 597553
rect 495438 597479 495494 597488
rect 498198 597544 498254 597553
rect 498198 597479 498254 597488
rect 500958 597544 501014 597553
rect 500958 597479 501014 597488
rect 452658 597408 452714 597417
rect 452658 597343 452714 597352
rect 452672 597038 452700 597343
rect 452660 597032 452712 597038
rect 452660 596974 452712 596980
rect 454038 597000 454094 597009
rect 454038 596935 454040 596944
rect 454092 596935 454094 596944
rect 455418 597000 455474 597009
rect 455418 596935 455474 596944
rect 454040 596906 454092 596912
rect 455432 596902 455460 596935
rect 455420 596896 455472 596902
rect 455420 596838 455472 596844
rect 449990 596456 450046 596465
rect 449990 596391 449992 596400
rect 450044 596391 450046 596400
rect 451094 596456 451150 596465
rect 451094 596391 451150 596400
rect 451278 596456 451334 596465
rect 451278 596391 451334 596400
rect 449992 596362 450044 596368
rect 451292 596358 451320 596391
rect 451280 596352 451332 596358
rect 451280 596294 451332 596300
rect 456798 596320 456854 596329
rect 456798 596255 456854 596264
rect 456812 596222 456840 596255
rect 456800 596216 456852 596222
rect 456800 596158 456852 596164
rect 462332 594425 462360 597479
rect 462318 594416 462374 594425
rect 462318 594351 462374 594360
rect 465092 594289 465120 597479
rect 465078 594280 465134 594289
rect 465078 594215 465134 594224
rect 467852 594153 467880 597479
rect 470598 596320 470654 596329
rect 470598 596255 470654 596264
rect 467838 594144 467894 594153
rect 467838 594079 467894 594088
rect 470612 594017 470640 596255
rect 470598 594008 470654 594017
rect 473372 593978 473400 597479
rect 474752 594046 474780 597479
rect 477512 594794 477540 597479
rect 480258 597000 480314 597009
rect 480258 596935 480314 596944
rect 477500 594788 477552 594794
rect 477500 594730 477552 594736
rect 480272 594726 480300 596935
rect 480260 594720 480312 594726
rect 480260 594662 480312 594668
rect 483032 594658 483060 597479
rect 483020 594652 483072 594658
rect 483020 594594 483072 594600
rect 485792 594590 485820 597479
rect 485780 594584 485832 594590
rect 485780 594526 485832 594532
rect 488552 594522 488580 597479
rect 492678 596728 492734 596737
rect 492678 596663 492734 596672
rect 489918 596320 489974 596329
rect 489918 596255 489974 596264
rect 488540 594516 488592 594522
rect 488540 594458 488592 594464
rect 489932 594454 489960 596255
rect 489920 594448 489972 594454
rect 489920 594390 489972 594396
rect 492692 594386 492720 596663
rect 492680 594380 492732 594386
rect 492680 594322 492732 594328
rect 495452 594318 495480 597479
rect 495440 594312 495492 594318
rect 495440 594254 495492 594260
rect 498212 594250 498240 597479
rect 498200 594244 498252 594250
rect 498200 594186 498252 594192
rect 500972 594182 501000 597479
rect 502338 597000 502394 597009
rect 502338 596935 502394 596944
rect 500960 594176 501012 594182
rect 500960 594118 501012 594124
rect 502352 594114 502380 596935
rect 505098 596864 505154 596873
rect 505098 596799 505154 596808
rect 502340 594108 502392 594114
rect 502340 594050 502392 594056
rect 474740 594040 474792 594046
rect 474740 593982 474792 593988
rect 470598 593943 470654 593952
rect 473360 593972 473412 593978
rect 473360 593914 473412 593920
rect 505112 592657 505140 596799
rect 505098 592648 505154 592657
rect 505098 592583 505154 592592
rect 449900 591320 449952 591326
rect 449900 591262 449952 591268
rect 536852 565894 536880 685850
rect 538218 679008 538274 679017
rect 538218 678943 538274 678952
rect 537484 643136 537536 643142
rect 537484 643078 537536 643084
rect 530952 565888 531004 565894
rect 530950 565856 530952 565865
rect 536840 565888 536892 565894
rect 531004 565856 531006 565865
rect 536840 565830 536892 565836
rect 530950 565791 531006 565800
rect 433338 563680 433394 563689
rect 433338 563615 433394 563624
rect 425520 478576 425572 478582
rect 425520 478518 425572 478524
rect 400128 477760 400180 477766
rect 400128 477702 400180 477708
rect 399944 477080 399996 477086
rect 399944 477022 399996 477028
rect 399852 476196 399904 476202
rect 399852 476138 399904 476144
rect 399760 476128 399812 476134
rect 399760 476070 399812 476076
rect 399956 470594 399984 477022
rect 400140 477018 400168 477702
rect 424140 477692 424192 477698
rect 424140 477634 424192 477640
rect 424152 477465 424180 477634
rect 425532 477465 425560 478518
rect 426624 478508 426676 478514
rect 426624 478450 426676 478456
rect 426164 477692 426216 477698
rect 426164 477634 426216 477640
rect 415398 477456 415454 477465
rect 415398 477391 415454 477400
rect 416778 477456 416834 477465
rect 416778 477391 416834 477400
rect 418158 477456 418214 477465
rect 418158 477391 418214 477400
rect 419538 477456 419594 477465
rect 419538 477391 419594 477400
rect 420918 477456 420974 477465
rect 420918 477391 420974 477400
rect 423126 477456 423182 477465
rect 423126 477391 423182 477400
rect 424138 477456 424194 477465
rect 424138 477391 424194 477400
rect 425518 477456 425574 477465
rect 425518 477391 425574 477400
rect 415412 477154 415440 477391
rect 416792 477222 416820 477391
rect 416780 477216 416832 477222
rect 416780 477158 416832 477164
rect 415400 477148 415452 477154
rect 415400 477090 415452 477096
rect 418172 477018 418200 477391
rect 419552 477086 419580 477391
rect 419540 477080 419592 477086
rect 419540 477022 419592 477028
rect 400128 477012 400180 477018
rect 400128 476954 400180 476960
rect 418160 477012 418212 477018
rect 418160 476954 418212 476960
rect 419540 476944 419592 476950
rect 419540 476886 419592 476892
rect 419552 476513 419580 476886
rect 420932 476814 420960 477391
rect 423140 476814 423168 477391
rect 420920 476808 420972 476814
rect 420920 476750 420972 476756
rect 423128 476808 423180 476814
rect 423128 476750 423180 476756
rect 425532 476746 425560 477391
rect 425520 476740 425572 476746
rect 425520 476682 425572 476688
rect 419538 476504 419594 476513
rect 426176 476474 426204 477634
rect 426636 477465 426664 478450
rect 427820 478440 427872 478446
rect 427820 478382 427872 478388
rect 428554 478408 428610 478417
rect 426622 477456 426678 477465
rect 426622 477391 426678 477400
rect 427726 477456 427782 477465
rect 427832 477442 427860 478382
rect 428554 478343 428610 478352
rect 430118 478408 430174 478417
rect 430118 478343 430120 478352
rect 428568 478310 428596 478343
rect 430172 478343 430174 478352
rect 430580 478372 430632 478378
rect 430120 478314 430172 478320
rect 430580 478314 430632 478320
rect 428556 478304 428608 478310
rect 428556 478246 428608 478252
rect 430028 478304 430080 478310
rect 430028 478246 430080 478252
rect 427782 477414 427860 477442
rect 427726 477391 427782 477400
rect 426636 477086 426664 477391
rect 427740 477154 427768 477391
rect 430040 477290 430068 478246
rect 430028 477284 430080 477290
rect 430028 477226 430080 477232
rect 430592 477222 430620 478314
rect 431314 478272 431370 478281
rect 431314 478207 431316 478216
rect 431368 478207 431370 478216
rect 432510 478272 432566 478281
rect 432510 478207 432566 478216
rect 433248 478236 433300 478242
rect 431316 478178 431368 478184
rect 432524 478174 432552 478207
rect 433248 478178 433300 478184
rect 432512 478168 432564 478174
rect 432512 478110 432564 478116
rect 433260 477426 433288 478178
rect 434628 478168 434680 478174
rect 434628 478110 434680 478116
rect 434444 477556 434496 477562
rect 434444 477498 434496 477504
rect 433432 477488 433484 477494
rect 433430 477456 433432 477465
rect 433484 477456 433486 477465
rect 433248 477420 433300 477426
rect 433430 477391 433486 477400
rect 433248 477362 433300 477368
rect 430580 477216 430632 477222
rect 430580 477158 430632 477164
rect 427728 477148 427780 477154
rect 427728 477090 427780 477096
rect 426624 477080 426676 477086
rect 426624 477022 426676 477028
rect 434456 476678 434484 477498
rect 434536 477488 434588 477494
rect 434534 477456 434536 477465
rect 434588 477456 434590 477465
rect 434534 477391 434590 477400
rect 434444 476672 434496 476678
rect 434444 476614 434496 476620
rect 433338 476504 433394 476513
rect 419538 476439 419594 476448
rect 426164 476468 426216 476474
rect 433338 476439 433394 476448
rect 426164 476410 426216 476416
rect 427818 476232 427874 476241
rect 427818 476167 427874 476176
rect 430578 476232 430634 476241
rect 430578 476167 430634 476176
rect 400128 476128 400180 476134
rect 400128 476070 400180 476076
rect 399680 470566 399984 470594
rect 399574 357096 399630 357105
rect 399574 357031 399630 357040
rect 399680 356969 399708 470566
rect 400140 444281 400168 476070
rect 427832 460193 427860 476167
rect 430592 461553 430620 476167
rect 433352 476134 433380 476439
rect 434640 476338 434668 478110
rect 436008 477624 436060 477630
rect 436008 477566 436060 477572
rect 435730 477456 435786 477465
rect 435730 477391 435786 477400
rect 435744 477018 435772 477391
rect 436020 477358 436048 477566
rect 436834 477456 436890 477465
rect 436834 477391 436890 477400
rect 438122 477456 438178 477465
rect 438122 477391 438178 477400
rect 442998 477456 443054 477465
rect 442998 477391 443054 477400
rect 447138 477456 447194 477465
rect 447138 477391 447194 477400
rect 448518 477456 448574 477465
rect 448518 477391 448520 477400
rect 436008 477352 436060 477358
rect 436008 477294 436060 477300
rect 435732 477012 435784 477018
rect 435732 476954 435784 476960
rect 435744 476406 435772 476954
rect 436848 476882 436876 477391
rect 438136 476950 438164 477391
rect 438858 477184 438914 477193
rect 438858 477119 438914 477128
rect 437480 476944 437532 476950
rect 437480 476886 437532 476892
rect 438124 476944 438176 476950
rect 438124 476886 438176 476892
rect 436836 476876 436888 476882
rect 436836 476818 436888 476824
rect 436848 476542 436876 476818
rect 437492 476610 437520 476886
rect 437480 476604 437532 476610
rect 437480 476546 437532 476552
rect 436836 476536 436888 476542
rect 436836 476478 436888 476484
rect 435732 476400 435784 476406
rect 435732 476342 435784 476348
rect 434628 476332 434680 476338
rect 434628 476274 434680 476280
rect 433340 476128 433392 476134
rect 433340 476070 433392 476076
rect 438872 473822 438900 477119
rect 440238 477048 440294 477057
rect 440238 476983 440294 476992
rect 438860 473816 438912 473822
rect 438860 473758 438912 473764
rect 440252 471986 440280 476983
rect 441618 476912 441674 476921
rect 441618 476847 441674 476856
rect 441632 476814 441660 476847
rect 441620 476808 441672 476814
rect 441620 476750 441672 476756
rect 443012 476746 443040 477391
rect 447152 477290 447180 477391
rect 448572 477391 448574 477400
rect 452658 477456 452714 477465
rect 452658 477391 452714 477400
rect 448520 477362 448572 477368
rect 452672 477358 452700 477391
rect 452660 477352 452712 477358
rect 452660 477294 452712 477300
rect 447140 477284 447192 477290
rect 447140 477226 447192 477232
rect 448520 477216 448572 477222
rect 444194 477184 444250 477193
rect 444194 477119 444250 477128
rect 444378 477184 444434 477193
rect 444378 477119 444434 477128
rect 445758 477184 445814 477193
rect 445758 477119 445760 477128
rect 444208 476814 444236 477119
rect 444392 477086 444420 477119
rect 445812 477119 445814 477128
rect 448518 477184 448520 477193
rect 448572 477184 448574 477193
rect 448518 477119 448574 477128
rect 451370 477184 451426 477193
rect 451370 477119 451426 477128
rect 458178 477184 458234 477193
rect 458178 477119 458234 477128
rect 462318 477184 462374 477193
rect 462318 477119 462374 477128
rect 445760 477090 445812 477096
rect 444380 477080 444432 477086
rect 445668 477080 445720 477086
rect 444380 477022 444432 477028
rect 445666 477048 445668 477057
rect 445720 477048 445722 477057
rect 445666 476983 445722 476992
rect 446402 477048 446458 477057
rect 446402 476983 446458 476992
rect 444196 476808 444248 476814
rect 444196 476750 444248 476756
rect 443000 476740 443052 476746
rect 443000 476682 443052 476688
rect 446416 476649 446444 476983
rect 451384 476678 451412 477119
rect 458192 477086 458220 477119
rect 458180 477080 458232 477086
rect 454038 477048 454094 477057
rect 454038 476983 454040 476992
rect 454092 476983 454094 476992
rect 456798 477048 456854 477057
rect 458180 477022 458232 477028
rect 456798 476983 456854 476992
rect 454040 476954 454092 476960
rect 456812 476950 456840 476983
rect 456800 476944 456852 476950
rect 455418 476912 455474 476921
rect 456800 476886 456852 476892
rect 456890 476912 456946 476921
rect 455418 476847 455420 476856
rect 455472 476847 455474 476856
rect 456890 476847 456946 476856
rect 455420 476818 455472 476824
rect 456904 476814 456932 476847
rect 456892 476808 456944 476814
rect 456892 476750 456944 476756
rect 451372 476672 451424 476678
rect 446402 476640 446458 476649
rect 451372 476614 451424 476620
rect 446402 476575 446458 476584
rect 441986 476504 442042 476513
rect 441986 476439 441988 476448
rect 442040 476439 442042 476448
rect 442998 476504 443054 476513
rect 442998 476439 443054 476448
rect 449898 476504 449954 476513
rect 449898 476439 449954 476448
rect 441988 476410 442040 476416
rect 443012 474609 443040 476439
rect 449912 476338 449940 476439
rect 449900 476332 449952 476338
rect 449900 476274 449952 476280
rect 445758 476232 445814 476241
rect 445758 476167 445814 476176
rect 447138 476232 447194 476241
rect 447138 476167 447194 476176
rect 449898 476232 449954 476241
rect 449898 476167 449954 476176
rect 442998 474600 443054 474609
rect 442998 474535 443054 474544
rect 440240 471980 440292 471986
rect 440240 471922 440292 471928
rect 445772 471510 445800 476167
rect 445760 471504 445812 471510
rect 445760 471446 445812 471452
rect 447152 471442 447180 476167
rect 447140 471436 447192 471442
rect 447140 471378 447192 471384
rect 449912 471374 449940 476167
rect 462332 474473 462360 477119
rect 483018 476912 483074 476921
rect 483018 476847 483074 476856
rect 474738 476504 474794 476513
rect 474738 476439 474794 476448
rect 477498 476504 477554 476513
rect 477498 476439 477554 476448
rect 465078 476232 465134 476241
rect 465078 476167 465134 476176
rect 467838 476232 467894 476241
rect 467838 476167 467894 476176
rect 470782 476232 470838 476241
rect 470782 476167 470838 476176
rect 473358 476232 473414 476241
rect 473358 476167 473414 476176
rect 462318 474464 462374 474473
rect 462318 474399 462374 474408
rect 465092 473890 465120 476167
rect 467852 474337 467880 476167
rect 467838 474328 467894 474337
rect 467838 474263 467894 474272
rect 470796 474201 470824 476167
rect 470782 474192 470838 474201
rect 470782 474127 470838 474136
rect 473372 474065 473400 476167
rect 473358 474056 473414 474065
rect 473358 473991 473414 474000
rect 474752 473958 474780 476439
rect 477512 474706 477540 476439
rect 480534 476232 480590 476241
rect 480534 476167 480590 476176
rect 477500 474700 477552 474706
rect 477500 474642 477552 474648
rect 480548 474638 480576 476167
rect 480536 474632 480588 474638
rect 480536 474574 480588 474580
rect 483032 474570 483060 476847
rect 490470 476776 490526 476785
rect 490470 476711 490526 476720
rect 498198 476776 498254 476785
rect 498198 476711 498254 476720
rect 485778 476232 485834 476241
rect 485778 476167 485834 476176
rect 488538 476232 488594 476241
rect 488538 476167 488594 476176
rect 483020 474564 483072 474570
rect 483020 474506 483072 474512
rect 485792 474502 485820 476167
rect 485780 474496 485832 474502
rect 485780 474438 485832 474444
rect 488552 474434 488580 476167
rect 488540 474428 488592 474434
rect 488540 474370 488592 474376
rect 490484 474366 490512 476711
rect 492678 476232 492734 476241
rect 492678 476167 492734 476176
rect 495438 476232 495494 476241
rect 495438 476167 495494 476176
rect 490472 474360 490524 474366
rect 490472 474302 490524 474308
rect 492692 474298 492720 476167
rect 492680 474292 492732 474298
rect 492680 474234 492732 474240
rect 495452 474162 495480 476167
rect 495440 474156 495492 474162
rect 495440 474098 495492 474104
rect 498212 474094 498240 476711
rect 502338 476368 502394 476377
rect 502338 476303 502394 476312
rect 500958 476232 501014 476241
rect 500958 476167 501014 476176
rect 498200 474088 498252 474094
rect 498200 474030 498252 474036
rect 500972 474026 501000 476167
rect 502352 474230 502380 476303
rect 505098 476232 505154 476241
rect 505098 476167 505154 476176
rect 502340 474224 502392 474230
rect 502340 474166 502392 474172
rect 500960 474020 501012 474026
rect 500960 473962 501012 473968
rect 474740 473952 474792 473958
rect 474740 473894 474792 473900
rect 465080 473884 465132 473890
rect 465080 473826 465132 473832
rect 449900 471368 449952 471374
rect 449900 471310 449952 471316
rect 505112 471306 505140 476167
rect 505100 471300 505152 471306
rect 505100 471242 505152 471248
rect 430578 461544 430634 461553
rect 430578 461479 430634 461488
rect 427818 460184 427874 460193
rect 427818 460119 427874 460128
rect 536852 447030 536880 565830
rect 530492 447024 530544 447030
rect 530492 446966 530544 446972
rect 536840 447024 536892 447030
rect 536840 446966 536892 446972
rect 530504 446457 530532 446966
rect 530490 446448 530546 446457
rect 530490 446383 530546 446392
rect 400126 444272 400182 444281
rect 400126 444207 400182 444216
rect 416042 358184 416098 358193
rect 416042 358119 416098 358128
rect 488538 358184 488594 358193
rect 488538 358119 488594 358128
rect 416056 358086 416084 358119
rect 416044 358080 416096 358086
rect 416044 358022 416096 358028
rect 423128 357400 423180 357406
rect 423126 357368 423128 357377
rect 423588 357400 423640 357406
rect 423180 357368 423182 357377
rect 423588 357342 423640 357348
rect 424966 357368 425022 357377
rect 423126 357303 423182 357312
rect 399666 356960 399722 356969
rect 399666 356895 399722 356904
rect 423600 356522 423628 357342
rect 424966 357303 425022 357312
rect 425426 357368 425482 357377
rect 425426 357303 425482 357312
rect 426898 357368 426954 357377
rect 426898 357303 426954 357312
rect 427634 357368 427690 357377
rect 427634 357303 427690 357312
rect 427818 357368 427874 357377
rect 427818 357303 427874 357312
rect 428554 357368 428610 357377
rect 428554 357303 428610 357312
rect 430026 357368 430082 357377
rect 430026 357303 430082 357312
rect 430578 357368 430634 357377
rect 430578 357303 430634 357312
rect 431958 357368 432014 357377
rect 431958 357303 432014 357312
rect 433338 357368 433394 357377
rect 434718 357368 434774 357377
rect 433338 357303 433394 357312
rect 433432 357332 433484 357338
rect 424980 356726 425008 357303
rect 424968 356720 425020 356726
rect 424968 356662 425020 356668
rect 423588 356516 423640 356522
rect 423588 356458 423640 356464
rect 424980 356250 425008 356662
rect 425440 356590 425468 357303
rect 426912 356658 426940 357303
rect 426900 356652 426952 356658
rect 426900 356594 426952 356600
rect 425428 356584 425480 356590
rect 425428 356526 425480 356532
rect 426348 356584 426400 356590
rect 426348 356526 426400 356532
rect 426360 356386 426388 356526
rect 426348 356380 426400 356386
rect 426348 356322 426400 356328
rect 426912 356318 426940 356594
rect 427648 356590 427676 357303
rect 427636 356584 427688 356590
rect 427636 356526 427688 356532
rect 426900 356312 426952 356318
rect 426900 356254 426952 356260
rect 424968 356244 425020 356250
rect 424968 356186 425020 356192
rect 399484 351076 399536 351082
rect 399484 351018 399536 351024
rect 427832 329118 427860 357303
rect 428568 356998 428596 357303
rect 428556 356992 428608 356998
rect 428556 356934 428608 356940
rect 428568 356658 428596 356934
rect 430040 356726 430068 357303
rect 429200 356720 429252 356726
rect 429200 356662 429252 356668
rect 430028 356720 430080 356726
rect 430028 356662 430080 356668
rect 428556 356652 428608 356658
rect 428556 356594 428608 356600
rect 429212 356454 429240 356662
rect 429200 356448 429252 356454
rect 429200 356390 429252 356396
rect 430592 330614 430620 357303
rect 430670 357232 430726 357241
rect 430670 357167 430726 357176
rect 430684 356930 430712 357167
rect 431972 357066 432000 357303
rect 431960 357060 432012 357066
rect 431960 357002 432012 357008
rect 430672 356924 430724 356930
rect 430672 356866 430724 356872
rect 430684 356454 430712 356866
rect 430672 356448 430724 356454
rect 430672 356390 430724 356396
rect 430580 330608 430632 330614
rect 430580 330550 430632 330556
rect 427820 329112 427872 329118
rect 427820 329054 427872 329060
rect 433352 297430 433380 357303
rect 434718 357303 434774 357312
rect 436834 357368 436890 357377
rect 436834 357303 436890 357312
rect 437478 357368 437534 357377
rect 437478 357303 437534 357312
rect 440238 357368 440294 357377
rect 440238 357303 440294 357312
rect 444286 357368 444342 357377
rect 444286 357303 444342 357312
rect 445850 357368 445906 357377
rect 445850 357303 445906 357312
rect 447230 357368 447286 357377
rect 447230 357303 447286 357312
rect 449898 357368 449954 357377
rect 449898 357303 449954 357312
rect 451462 357368 451518 357377
rect 451462 357303 451518 357312
rect 452658 357368 452714 357377
rect 452658 357303 452714 357312
rect 454682 357368 454738 357377
rect 454682 357303 454738 357312
rect 457534 357368 457590 357377
rect 457534 357303 457590 357312
rect 462318 357368 462374 357377
rect 462318 357303 462374 357312
rect 464342 357368 464398 357377
rect 464342 357303 464398 357312
rect 467838 357368 467894 357377
rect 467838 357303 467894 357312
rect 472622 357368 472678 357377
rect 472622 357303 472678 357312
rect 477498 357368 477554 357377
rect 477498 357303 477554 357312
rect 485778 357368 485834 357377
rect 485778 357303 485834 357312
rect 433432 357274 433484 357280
rect 433444 357241 433472 357274
rect 433430 357232 433486 357241
rect 433430 357167 433486 357176
rect 434626 357232 434682 357241
rect 434626 357167 434628 357176
rect 434680 357167 434682 357176
rect 434628 357138 434680 357144
rect 434640 356930 434668 357138
rect 434628 356924 434680 356930
rect 434628 356866 434680 356872
rect 434732 331906 434760 357303
rect 436006 357232 436062 357241
rect 436006 357167 436062 357176
rect 436020 357134 436048 357167
rect 436008 357128 436060 357134
rect 436008 357070 436060 357076
rect 436020 356998 436048 357070
rect 436008 356992 436060 356998
rect 436008 356934 436060 356940
rect 436848 356862 436876 357303
rect 436836 356856 436888 356862
rect 436836 356798 436888 356804
rect 436848 356182 436876 356798
rect 436836 356176 436888 356182
rect 436836 356118 436888 356124
rect 437492 342922 437520 357303
rect 438398 357232 438454 357241
rect 438398 357167 438454 357176
rect 438412 356794 438440 357167
rect 437572 356788 437624 356794
rect 437572 356730 437624 356736
rect 438400 356788 438452 356794
rect 438400 356730 438452 356736
rect 437584 356114 437612 356730
rect 437572 356108 437624 356114
rect 437572 356050 437624 356056
rect 437480 342916 437532 342922
rect 437480 342858 437532 342864
rect 434720 331900 434772 331906
rect 434720 331842 434772 331848
rect 440252 327826 440280 357303
rect 444300 357270 444328 357303
rect 444288 357264 444340 357270
rect 443090 357232 443146 357241
rect 444288 357206 444340 357212
rect 443090 357167 443146 357176
rect 441710 356552 441766 356561
rect 441710 356487 441712 356496
rect 441764 356487 441766 356496
rect 442998 356552 443054 356561
rect 442998 356487 443054 356496
rect 441712 356458 441764 356464
rect 441986 356416 442042 356425
rect 443012 356386 443040 356487
rect 441986 356351 442042 356360
rect 443000 356380 443052 356386
rect 442000 356250 442028 356351
rect 443000 356322 443052 356328
rect 441988 356244 442040 356250
rect 441988 356186 442040 356192
rect 443104 341630 443132 357167
rect 445668 357128 445720 357134
rect 445666 357096 445668 357105
rect 445720 357096 445722 357105
rect 445666 357031 445722 357040
rect 445758 356688 445814 356697
rect 445758 356623 445814 356632
rect 445772 356590 445800 356623
rect 445760 356584 445812 356590
rect 445760 356526 445812 356532
rect 444378 356416 444434 356425
rect 444378 356351 444434 356360
rect 444392 356318 444420 356351
rect 444380 356312 444432 356318
rect 444380 356254 444432 356260
rect 443092 341624 443144 341630
rect 443092 341566 443144 341572
rect 445864 336054 445892 357303
rect 447138 357096 447194 357105
rect 447138 357031 447194 357040
rect 447152 356658 447180 357031
rect 447140 356652 447192 356658
rect 447140 356594 447192 356600
rect 447244 344418 447272 357303
rect 448518 356824 448574 356833
rect 448518 356759 448574 356768
rect 448532 356726 448560 356759
rect 448520 356720 448572 356726
rect 448520 356662 448572 356668
rect 448518 356552 448574 356561
rect 448518 356487 448574 356496
rect 448532 356454 448560 356487
rect 448520 356448 448572 356454
rect 448520 356390 448572 356396
rect 449912 349858 449940 357303
rect 451476 357202 451504 357303
rect 451464 357196 451516 357202
rect 451464 357138 451516 357144
rect 449990 357096 450046 357105
rect 449990 357031 449992 357040
rect 450044 357031 450046 357040
rect 449992 357002 450044 357008
rect 449900 349852 449952 349858
rect 449900 349794 449952 349800
rect 447232 344412 447284 344418
rect 447232 344354 447284 344360
rect 452672 337414 452700 357303
rect 454038 357096 454094 357105
rect 454038 357031 454094 357040
rect 454052 356998 454080 357031
rect 454040 356992 454092 356998
rect 452750 356960 452806 356969
rect 454040 356934 454092 356940
rect 452750 356895 452752 356904
rect 452804 356895 452806 356904
rect 452752 356866 452804 356872
rect 452660 337408 452712 337414
rect 452660 337350 452712 337356
rect 445852 336048 445904 336054
rect 445852 335990 445904 335996
rect 440240 327820 440292 327826
rect 440240 327762 440292 327768
rect 454696 305658 454724 357303
rect 456800 357264 456852 357270
rect 456798 357232 456800 357241
rect 456852 357232 456854 357241
rect 456798 357167 456854 357176
rect 455418 356960 455474 356969
rect 455418 356895 455474 356904
rect 455432 356862 455460 356895
rect 455420 356856 455472 356862
rect 455420 356798 455472 356804
rect 456798 356824 456854 356833
rect 456798 356759 456800 356768
rect 456852 356759 456854 356768
rect 456800 356730 456852 356736
rect 457444 356108 457496 356114
rect 457444 356050 457496 356056
rect 454684 305652 454736 305658
rect 454684 305594 454736 305600
rect 457456 304298 457484 356050
rect 457548 320958 457576 357303
rect 458178 357232 458234 357241
rect 458178 357167 458234 357176
rect 458192 357134 458220 357167
rect 458180 357128 458232 357134
rect 458180 357070 458232 357076
rect 460938 356144 460994 356153
rect 460938 356079 460940 356088
rect 460992 356079 460994 356088
rect 460940 356050 460992 356056
rect 457536 320952 457588 320958
rect 457536 320894 457588 320900
rect 457444 304292 457496 304298
rect 457444 304234 457496 304240
rect 433340 297424 433392 297430
rect 433340 297366 433392 297372
rect 462332 293282 462360 357303
rect 464356 316742 464384 357303
rect 467852 356658 467880 357303
rect 464436 356652 464488 356658
rect 464436 356594 464488 356600
rect 467840 356652 467892 356658
rect 467840 356594 467892 356600
rect 464448 318102 464476 356594
rect 471244 356516 471296 356522
rect 471244 356458 471296 356464
rect 467196 356312 467248 356318
rect 467196 356254 467248 356260
rect 470782 356280 470838 356289
rect 467104 356108 467156 356114
rect 467104 356050 467156 356056
rect 464436 318096 464488 318102
rect 464436 318038 464488 318044
rect 464344 316736 464396 316742
rect 464344 316678 464396 316684
rect 467116 300150 467144 356050
rect 467208 308446 467236 356254
rect 470782 356215 470838 356224
rect 470796 356114 470824 356215
rect 470784 356108 470836 356114
rect 470784 356050 470836 356056
rect 467196 308440 467248 308446
rect 467196 308382 467248 308388
rect 471256 307086 471284 356458
rect 471244 307080 471296 307086
rect 471244 307022 471296 307028
rect 472636 301510 472664 357303
rect 477512 356522 477540 357303
rect 480534 357096 480590 357105
rect 480534 357031 480590 357040
rect 477500 356516 477552 356522
rect 477500 356458 477552 356464
rect 474738 356416 474794 356425
rect 474738 356351 474794 356360
rect 479524 356380 479576 356386
rect 474752 356318 474780 356351
rect 479524 356322 479576 356328
rect 474740 356312 474792 356318
rect 474740 356254 474792 356260
rect 476764 356312 476816 356318
rect 476764 356254 476816 356260
rect 472716 356176 472768 356182
rect 472716 356118 472768 356124
rect 472728 315382 472756 356118
rect 472716 315376 472768 315382
rect 472716 315318 472768 315324
rect 476776 302938 476804 356254
rect 476856 356108 476908 356114
rect 476856 356050 476908 356056
rect 476868 311166 476896 356050
rect 476856 311160 476908 311166
rect 476856 311102 476908 311108
rect 476764 302932 476816 302938
rect 476764 302874 476816 302880
rect 472624 301504 472676 301510
rect 472624 301446 472676 301452
rect 467104 300144 467156 300150
rect 467104 300086 467156 300092
rect 479536 297498 479564 356322
rect 480548 356182 480576 357031
rect 483018 356552 483074 356561
rect 483018 356487 483074 356496
rect 483032 356318 483060 356487
rect 483020 356312 483072 356318
rect 483020 356254 483072 356260
rect 482284 356244 482336 356250
rect 482284 356186 482336 356192
rect 480536 356176 480588 356182
rect 480536 356118 480588 356124
rect 479524 297492 479576 297498
rect 479524 297434 479576 297440
rect 482296 296002 482324 356186
rect 482284 295996 482336 296002
rect 482284 295938 482336 295944
rect 462320 293276 462372 293282
rect 462320 293218 462372 293224
rect 485792 291854 485820 357303
rect 488552 356386 488580 358119
rect 498198 357368 498254 357377
rect 498198 357303 498254 357312
rect 498212 356930 498240 357303
rect 491944 356924 491996 356930
rect 491944 356866 491996 356872
rect 498200 356924 498252 356930
rect 498200 356866 498252 356872
rect 488540 356380 488592 356386
rect 488540 356322 488592 356328
rect 489918 356280 489974 356289
rect 489918 356215 489920 356224
rect 489972 356215 489974 356224
rect 489920 356186 489972 356192
rect 487804 356176 487856 356182
rect 487804 356118 487856 356124
rect 487816 309806 487844 356118
rect 491956 319530 491984 356866
rect 502338 356824 502394 356833
rect 502338 356759 502394 356768
rect 500958 356416 501014 356425
rect 500958 356351 501014 356360
rect 500972 356318 501000 356351
rect 494704 356312 494756 356318
rect 500960 356312 501012 356318
rect 494704 356254 494756 356260
rect 495438 356280 495494 356289
rect 492678 356144 492734 356153
rect 492678 356079 492680 356088
rect 492732 356079 492734 356088
rect 492680 356050 492732 356056
rect 491944 319524 491996 319530
rect 491944 319466 491996 319472
rect 494716 313954 494744 356254
rect 500960 356254 501012 356260
rect 495438 356215 495494 356224
rect 495452 356182 495480 356215
rect 495440 356176 495492 356182
rect 495440 356118 495492 356124
rect 497464 356108 497516 356114
rect 497464 356050 497516 356056
rect 494704 313948 494756 313954
rect 494704 313890 494756 313896
rect 487804 309800 487856 309806
rect 487804 309742 487856 309748
rect 497476 294642 497504 356050
rect 497464 294636 497516 294642
rect 497464 294578 497516 294584
rect 485780 291848 485832 291854
rect 485780 291790 485832 291796
rect 502352 290494 502380 356759
rect 505098 356144 505154 356153
rect 505098 356079 505100 356088
rect 505152 356079 505154 356088
rect 505100 356050 505152 356056
rect 537496 322250 537524 643078
rect 537668 563100 537720 563106
rect 537668 563042 537720 563048
rect 537576 510672 537628 510678
rect 537576 510614 537628 510620
rect 537484 322244 537536 322250
rect 537484 322186 537536 322192
rect 502340 290488 502392 290494
rect 502340 290430 502392 290436
rect 396724 289808 396776 289814
rect 396724 289750 396776 289756
rect 449900 287496 449952 287502
rect 449900 287438 449952 287444
rect 364340 286476 364392 286482
rect 364340 286418 364392 286424
rect 361672 279812 361724 279818
rect 361672 279754 361724 279760
rect 361684 248414 361712 279754
rect 364352 248414 364380 286418
rect 368480 286408 368532 286414
rect 368480 286350 368532 286356
rect 367100 280628 367152 280634
rect 367100 280570 367152 280576
rect 361684 248386 362264 248414
rect 364352 248386 364656 248414
rect 362236 229922 362264 248386
rect 364628 229922 364656 248386
rect 367112 229922 367140 280570
rect 368492 248414 368520 286350
rect 374000 286340 374052 286346
rect 374000 286282 374052 286288
rect 371240 285116 371292 285122
rect 371240 285058 371292 285064
rect 371252 248414 371280 285058
rect 374012 248414 374040 286282
rect 378140 286272 378192 286278
rect 378140 286214 378192 286220
rect 376760 285048 376812 285054
rect 376760 284990 376812 284996
rect 368492 248386 369440 248414
rect 371252 248386 371832 248414
rect 374012 248386 374224 248414
rect 369412 229922 369440 248386
rect 371804 229922 371832 248386
rect 374196 229922 374224 248386
rect 376772 229922 376800 284990
rect 378152 248414 378180 286214
rect 383660 286204 383712 286210
rect 383660 286146 383712 286152
rect 380900 283756 380952 283762
rect 380900 283698 380952 283704
rect 380912 248414 380940 283698
rect 383672 248414 383700 286146
rect 387800 286136 387852 286142
rect 387800 286078 387852 286084
rect 386420 284980 386472 284986
rect 386420 284922 386472 284928
rect 378152 248386 379008 248414
rect 380912 248386 381400 248414
rect 383672 248386 383792 248414
rect 378980 229922 379008 248386
rect 381372 229922 381400 248386
rect 383764 229922 383792 248386
rect 386432 229922 386460 284922
rect 387812 248414 387840 286078
rect 402980 286068 403032 286074
rect 402980 286010 403032 286016
rect 396080 284912 396132 284918
rect 396080 284854 396132 284860
rect 393320 283688 393372 283694
rect 393320 283630 393372 283636
rect 390560 279676 390612 279682
rect 390560 279618 390612 279624
rect 390572 248414 390600 279618
rect 387812 248386 388576 248414
rect 390572 248386 390968 248414
rect 388548 229922 388576 248386
rect 390940 229922 390968 248386
rect 393332 229922 393360 283630
rect 362236 229894 362618 229922
rect 364628 229894 365010 229922
rect 367112 229894 367402 229922
rect 369412 229894 369794 229922
rect 371804 229894 372186 229922
rect 374196 229894 374578 229922
rect 376772 229894 376970 229922
rect 378980 229894 379362 229922
rect 381372 229894 381754 229922
rect 383764 229894 384146 229922
rect 386432 229894 386538 229922
rect 388548 229894 388930 229922
rect 390940 229894 391322 229922
rect 393332 229894 393714 229922
rect 396092 229908 396120 284854
rect 397460 284844 397512 284850
rect 397460 284786 397512 284792
rect 397472 248414 397500 284786
rect 400220 280560 400272 280566
rect 400220 280502 400272 280508
rect 400232 248414 400260 280502
rect 397472 248386 398144 248414
rect 400232 248386 400536 248414
rect 398116 229922 398144 248386
rect 400508 229922 400536 248386
rect 402992 229922 403020 286010
rect 404360 286000 404412 286006
rect 404360 285942 404412 285948
rect 404372 248414 404400 285942
rect 407120 285932 407172 285938
rect 407120 285874 407172 285880
rect 407132 248414 407160 285874
rect 412640 285864 412692 285870
rect 412640 285806 412692 285812
rect 409880 279608 409932 279614
rect 409880 279550 409932 279556
rect 409892 248414 409920 279550
rect 404372 248386 405320 248414
rect 407132 248386 407712 248414
rect 409892 248386 410104 248414
rect 405292 229922 405320 248386
rect 407684 229922 407712 248386
rect 410076 229922 410104 248386
rect 412652 229922 412680 285806
rect 416780 285796 416832 285802
rect 416780 285738 416832 285744
rect 414020 284776 414072 284782
rect 414020 284718 414072 284724
rect 414032 248414 414060 284718
rect 416792 248414 416820 285738
rect 422300 285728 422352 285734
rect 422300 285670 422352 285676
rect 419540 284708 419592 284714
rect 419540 284650 419592 284656
rect 419552 248414 419580 284650
rect 414032 248386 414888 248414
rect 416792 248386 417280 248414
rect 419552 248386 419672 248414
rect 414860 229922 414888 248386
rect 417252 229922 417280 248386
rect 419644 229922 419672 248386
rect 422312 229922 422340 285670
rect 423680 284640 423732 284646
rect 423680 284582 423732 284588
rect 423692 248414 423720 284582
rect 426440 284572 426492 284578
rect 426440 284514 426492 284520
rect 426452 248414 426480 284514
rect 429200 284504 429252 284510
rect 429200 284446 429252 284452
rect 423692 248386 424456 248414
rect 426452 248386 426848 248414
rect 424428 229922 424456 248386
rect 426820 229922 426848 248386
rect 429212 229922 429240 284446
rect 436100 284436 436152 284442
rect 436100 284378 436152 284384
rect 433340 283552 433392 283558
rect 433340 283494 433392 283500
rect 431960 280968 432012 280974
rect 431960 280910 432012 280916
rect 398116 229894 398498 229922
rect 400508 229894 400890 229922
rect 402992 229894 403282 229922
rect 405292 229894 405674 229922
rect 407684 229894 408066 229922
rect 410076 229894 410458 229922
rect 412652 229894 412850 229922
rect 414860 229894 415242 229922
rect 417252 229894 417634 229922
rect 419644 229894 420026 229922
rect 422312 229894 422418 229922
rect 424428 229894 424810 229922
rect 426820 229894 427202 229922
rect 429212 229894 429594 229922
rect 431972 229908 432000 280910
rect 433352 248414 433380 283494
rect 436112 248414 436140 284378
rect 448520 284368 448572 284374
rect 448520 284310 448572 284316
rect 440240 280492 440292 280498
rect 440240 280434 440292 280440
rect 438860 280424 438912 280430
rect 438860 280366 438912 280372
rect 433352 248386 434024 248414
rect 436112 248386 436416 248414
rect 433996 229922 434024 248386
rect 436388 229922 436416 248386
rect 438872 229922 438900 280366
rect 440252 248414 440280 280434
rect 443000 280356 443052 280362
rect 443000 280298 443052 280304
rect 443012 248414 443040 280298
rect 445760 280288 445812 280294
rect 445760 280230 445812 280236
rect 445772 248414 445800 280230
rect 440252 248386 441200 248414
rect 443012 248386 443592 248414
rect 445772 248386 445984 248414
rect 441172 229922 441200 248386
rect 443564 229922 443592 248386
rect 445956 229922 445984 248386
rect 448532 229922 448560 284310
rect 449912 248414 449940 287438
rect 458180 287428 458232 287434
rect 458180 287370 458232 287376
rect 456062 282024 456118 282033
rect 456062 281959 456118 281968
rect 453304 281716 453356 281722
rect 453304 281658 453356 281664
rect 449912 248386 450768 248414
rect 450740 229922 450768 248386
rect 453316 233034 453344 281658
rect 453212 233028 453264 233034
rect 453212 232970 453264 232976
rect 453304 233028 453356 233034
rect 453304 232970 453356 232976
rect 453224 229922 453252 232970
rect 456076 232966 456104 281959
rect 455880 232960 455932 232966
rect 455880 232902 455932 232908
rect 456064 232960 456116 232966
rect 456064 232902 456116 232908
rect 433996 229894 434378 229922
rect 436388 229894 436770 229922
rect 438872 229894 439162 229922
rect 441172 229894 441554 229922
rect 443564 229894 443946 229922
rect 445956 229894 446338 229922
rect 448532 229894 448730 229922
rect 450740 229894 451122 229922
rect 453224 229894 453514 229922
rect 455892 229908 455920 232902
rect 458192 229922 458220 287370
rect 471980 287360 472032 287366
rect 471980 287302 472032 287308
rect 469862 281888 469918 281897
rect 469862 281823 469918 281832
rect 459560 281784 459612 281790
rect 459560 281726 459612 281732
rect 459572 248414 459600 281726
rect 462320 281648 462372 281654
rect 462320 281590 462372 281596
rect 462332 248414 462360 281590
rect 467840 279744 467892 279750
rect 467840 279686 467892 279692
rect 459572 248386 460336 248414
rect 462332 248386 462728 248414
rect 460308 229922 460336 248386
rect 462700 229922 462728 248386
rect 465448 233980 465500 233986
rect 465448 233922 465500 233928
rect 458192 229894 458298 229922
rect 460308 229894 460690 229922
rect 462700 229894 463082 229922
rect 465460 229908 465488 233922
rect 467852 229908 467880 279686
rect 469876 232898 469904 281823
rect 471992 248414 472020 287302
rect 474740 287292 474792 287298
rect 474740 287234 474792 287240
rect 471992 248386 472296 248414
rect 469772 232892 469824 232898
rect 469772 232834 469824 232840
rect 469864 232892 469916 232898
rect 469864 232834 469916 232840
rect 469784 229922 469812 232834
rect 472268 229922 472296 248386
rect 474752 229922 474780 287234
rect 478880 287224 478932 287230
rect 478880 287166 478932 287172
rect 517518 287192 517574 287201
rect 476120 280900 476172 280906
rect 476120 280842 476172 280848
rect 476132 248414 476160 280842
rect 478892 248414 478920 287166
rect 484400 287156 484452 287162
rect 517518 287127 517574 287136
rect 484400 287098 484452 287104
rect 481640 281580 481692 281586
rect 481640 281522 481692 281528
rect 481652 248414 481680 281522
rect 476132 248386 477080 248414
rect 478892 248386 479472 248414
rect 481652 248386 481864 248414
rect 477052 229922 477080 248386
rect 479444 229922 479472 248386
rect 481836 229922 481864 248386
rect 484412 229922 484440 287098
rect 485780 287088 485832 287094
rect 485780 287030 485832 287036
rect 485792 248414 485820 287030
rect 491942 281752 491998 281761
rect 491942 281687 491998 281696
rect 491300 279880 491352 279886
rect 491300 279822 491352 279828
rect 491312 248414 491340 279822
rect 485792 248386 486648 248414
rect 491312 248386 491432 248414
rect 486620 229922 486648 248386
rect 489368 233028 489420 233034
rect 489368 232970 489420 232976
rect 469784 229894 470258 229922
rect 472268 229894 472650 229922
rect 474752 229894 475042 229922
rect 477052 229894 477434 229922
rect 479444 229894 479826 229922
rect 481836 229894 482218 229922
rect 484412 229894 484610 229922
rect 486620 229894 487002 229922
rect 489380 229908 489408 232970
rect 491404 229922 491432 248386
rect 491956 233034 491984 281687
rect 514758 281616 514814 281625
rect 514758 281551 514814 281560
rect 511264 280220 511316 280226
rect 511264 280162 511316 280168
rect 505100 279540 505152 279546
rect 505100 279482 505152 279488
rect 505112 248414 505140 279482
rect 505112 248386 505784 248414
rect 494152 233912 494204 233918
rect 494152 233854 494204 233860
rect 498934 233880 498990 233889
rect 491944 233028 491996 233034
rect 491944 232970 491996 232976
rect 491404 229894 491786 229922
rect 494164 229908 494192 233854
rect 498934 233815 498990 233824
rect 496544 232824 496596 232830
rect 496544 232766 496596 232772
rect 496556 229908 496584 232766
rect 498948 229908 498976 233815
rect 503720 233028 503772 233034
rect 503720 232970 503772 232976
rect 501328 232756 501380 232762
rect 501328 232698 501380 232704
rect 501340 229908 501368 232698
rect 503732 229908 503760 232970
rect 505756 229922 505784 248386
rect 508504 232688 508556 232694
rect 508504 232630 508556 232636
rect 505756 229894 506138 229922
rect 508516 229908 508544 232630
rect 511276 232626 511304 280162
rect 514772 248414 514800 281551
rect 517532 248414 517560 287127
rect 537588 283626 537616 510614
rect 537680 344350 537708 563042
rect 538232 559201 538260 678943
rect 538864 670744 538916 670750
rect 538864 670686 538916 670692
rect 538218 559192 538274 559201
rect 538218 559127 538274 559136
rect 538232 454782 538260 559127
rect 538220 454776 538272 454782
rect 538220 454718 538272 454724
rect 538232 439793 538260 454718
rect 538218 439784 538274 439793
rect 538218 439719 538274 439728
rect 537668 344344 537720 344350
rect 537668 344286 537720 344292
rect 538876 340202 538904 670686
rect 538956 616888 539008 616894
rect 538956 616830 539008 616836
rect 538864 340196 538916 340202
rect 538864 340138 538916 340144
rect 538968 326398 538996 616830
rect 541624 524476 541676 524482
rect 541624 524418 541676 524424
rect 540244 484424 540296 484430
rect 540244 484366 540296 484372
rect 538956 326392 539008 326398
rect 538956 326334 539008 326340
rect 540256 320890 540284 484366
rect 540336 404388 540388 404394
rect 540336 404330 540388 404336
rect 540348 347070 540376 404330
rect 540336 347064 540388 347070
rect 540336 347006 540388 347012
rect 540244 320884 540296 320890
rect 540244 320826 540296 320832
rect 541636 315314 541664 524418
rect 541624 315308 541676 315314
rect 541624 315250 541676 315256
rect 542372 290601 542400 702406
rect 544384 536852 544436 536858
rect 544384 536794 544436 536800
rect 543004 364404 543056 364410
rect 543004 364346 543056 364352
rect 543016 327758 543044 364346
rect 543004 327752 543056 327758
rect 543004 327694 543056 327700
rect 542358 290592 542414 290601
rect 542358 290527 542414 290536
rect 544396 284889 544424 536794
rect 548524 430636 548576 430642
rect 548524 430578 548576 430584
rect 547144 378208 547196 378214
rect 547144 378150 547196 378156
rect 547156 289134 547184 378150
rect 548536 290465 548564 430578
rect 558932 345710 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 558920 345704 558972 345710
rect 558920 345646 558972 345652
rect 580276 338774 580304 683839
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580368 353977 580396 630799
rect 580446 418296 580502 418305
rect 580446 418231 580502 418240
rect 580354 353968 580410 353977
rect 580354 353903 580410 353912
rect 580460 348430 580488 418231
rect 580448 348424 580500 348430
rect 580448 348366 580500 348372
rect 580264 338768 580316 338774
rect 580264 338710 580316 338716
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 548522 290456 548578 290465
rect 548522 290391 548578 290400
rect 547144 289128 547196 289134
rect 547144 289070 547196 289076
rect 544382 284880 544438 284889
rect 544382 284815 544438 284824
rect 537576 283620 537628 283626
rect 537576 283562 537628 283568
rect 580540 283484 580592 283490
rect 580540 283426 580592 283432
rect 538956 283348 539008 283354
rect 538956 283290 539008 283296
rect 538864 283212 538916 283218
rect 538864 283154 538916 283160
rect 514772 248386 515352 248414
rect 517532 248386 517744 248414
rect 510896 232620 510948 232626
rect 510896 232562 510948 232568
rect 511264 232620 511316 232626
rect 511264 232562 511316 232568
rect 510908 229908 510936 232562
rect 513286 232520 513342 232529
rect 513286 232455 513342 232464
rect 513300 229908 513328 232455
rect 515324 229922 515352 248386
rect 517716 229922 517744 248386
rect 520464 232960 520516 232966
rect 520464 232902 520516 232908
rect 515324 229894 515706 229922
rect 517716 229894 518098 229922
rect 520476 229908 520504 232902
rect 525248 232892 525300 232898
rect 525248 232834 525300 232840
rect 522856 232552 522908 232558
rect 522856 232494 522908 232500
rect 522868 229908 522896 232494
rect 525260 229908 525288 232834
rect 527640 232620 527692 232626
rect 527640 232562 527692 232568
rect 527652 229908 527680 232562
rect 537208 231872 537260 231878
rect 537208 231814 537260 231820
rect 534814 230616 534870 230625
rect 534814 230551 534870 230560
rect 530032 230512 530084 230518
rect 530032 230454 530084 230460
rect 530044 229908 530072 230454
rect 534828 229908 534856 230551
rect 537220 229908 537248 231814
rect 532413 229200 532422 229256
rect 532478 229200 532487 229256
rect 538876 84194 538904 283154
rect 538968 86970 538996 283290
rect 540244 283280 540296 283286
rect 540244 283222 540296 283228
rect 540256 126954 540284 283222
rect 543096 283144 543148 283150
rect 543096 283086 543148 283092
rect 543004 283008 543056 283014
rect 543004 282950 543056 282956
rect 540334 280256 540390 280265
rect 540334 280191 540390 280200
rect 540348 139398 540376 280191
rect 540336 139392 540388 139398
rect 540336 139334 540388 139340
rect 540244 126948 540296 126954
rect 540244 126890 540296 126896
rect 543016 113150 543044 282950
rect 543108 167006 543136 283086
rect 544384 283076 544436 283082
rect 544384 283018 544436 283024
rect 544396 206990 544424 283018
rect 580356 282940 580408 282946
rect 580356 282882 580408 282888
rect 580262 280936 580318 280945
rect 580262 280871 580318 280880
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 544384 206984 544436 206990
rect 544384 206926 544436 206932
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 543096 167000 543148 167006
rect 543096 166942 543148 166948
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 139392 579856 139398
rect 579802 139360 579804 139369
rect 579856 139360 579858 139369
rect 579802 139295 579858 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 543004 113144 543056 113150
rect 543004 113086 543056 113092
rect 579620 113144 579672 113150
rect 579620 113086 579672 113092
rect 579632 112849 579660 113086
rect 579618 112840 579674 112849
rect 579618 112775 579674 112784
rect 538956 86964 539008 86970
rect 538956 86906 539008 86912
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 538876 84166 538996 84194
rect 538968 73166 538996 84166
rect 538956 73160 539008 73166
rect 538956 73102 539008 73108
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580276 59673 580304 280871
rect 580368 152697 580396 282882
rect 580446 280800 580502 280809
rect 580446 280735 580502 280744
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 580460 99521 580488 280735
rect 580552 179217 580580 283426
rect 580724 283416 580776 283422
rect 580724 283358 580776 283364
rect 580632 280832 580684 280838
rect 580632 280774 580684 280780
rect 580644 192545 580672 280774
rect 580736 219065 580764 283358
rect 580722 219056 580778 219065
rect 580722 218991 580778 219000
rect 580630 192536 580686 192545
rect 580630 192471 580686 192480
rect 580538 179208 580594 179217
rect 580538 179143 580594 179152
rect 580446 99512 580502 99521
rect 580446 99447 580502 99456
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 367100 49020 367152 49026
rect 367100 48962 367152 48968
rect 361580 48204 361632 48210
rect 361580 48146 361632 48152
rect 346400 44940 346452 44946
rect 346400 44882 346452 44888
rect 346412 16574 346440 44882
rect 353300 36576 353352 36582
rect 353300 36518 353352 36524
rect 349160 19984 349212 19990
rect 349160 19926 349212 19932
rect 346412 16546 346992 16574
rect 332692 6384 332744 6390
rect 332692 6326 332744 6332
rect 331864 3528 331916 3534
rect 331864 3470 331916 3476
rect 332704 480 332732 6326
rect 336280 6316 336332 6322
rect 336280 6258 336332 6264
rect 336292 480 336320 6258
rect 339868 6248 339920 6254
rect 339868 6190 339920 6196
rect 339880 480 339908 6190
rect 343364 6180 343416 6186
rect 343364 6122 343416 6128
rect 343376 480 343404 6122
rect 346964 480 346992 16546
rect 349172 2378 349200 19926
rect 353312 16574 353340 36518
rect 357440 35216 357492 35222
rect 357440 35158 357492 35164
rect 357452 16574 357480 35158
rect 364340 21480 364392 21486
rect 364340 21422 364392 21428
rect 360200 18692 360252 18698
rect 360200 18634 360252 18640
rect 360212 16574 360240 18634
rect 364352 16574 364380 21422
rect 367112 16574 367140 48962
rect 404924 48210 404952 50116
rect 494900 48278 494928 50116
rect 494888 48272 494940 48278
rect 494888 48214 494940 48220
rect 404912 48204 404964 48210
rect 404912 48146 404964 48152
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 416780 44872 416832 44878
rect 416780 44814 416832 44820
rect 385040 43512 385092 43518
rect 385040 43454 385092 43460
rect 371240 38004 371292 38010
rect 371240 37946 371292 37952
rect 353312 16546 353616 16574
rect 357452 16546 357572 16574
rect 360212 16546 361160 16574
rect 364352 16546 364656 16574
rect 367112 16546 367784 16574
rect 349160 2372 349212 2378
rect 349160 2314 349212 2320
rect 350448 2372 350500 2378
rect 350448 2314 350500 2320
rect 350460 480 350488 2314
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 357544 480 357572 16546
rect 361132 480 361160 16546
rect 364628 480 364656 16546
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 37946
rect 382280 29708 382332 29714
rect 382280 29650 382332 29656
rect 378140 26988 378192 26994
rect 378140 26930 378192 26936
rect 374000 25628 374052 25634
rect 374000 25570 374052 25576
rect 374012 3398 374040 25570
rect 378152 16574 378180 26930
rect 382292 16574 382320 29650
rect 385052 16574 385080 43454
rect 396080 39432 396132 39438
rect 396080 39374 396132 39380
rect 391940 33788 391992 33794
rect 391940 33730 391992 33736
rect 389180 31068 389232 31074
rect 389180 31010 389232 31016
rect 389192 16574 389220 31010
rect 391952 16574 391980 33730
rect 378152 16546 378456 16574
rect 382292 16546 382412 16574
rect 385052 16546 386000 16574
rect 389192 16546 389496 16574
rect 391952 16546 392624 16574
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 382384 480 382412 16546
rect 385972 480 386000 16546
rect 389468 480 389496 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 39374
rect 414020 28348 414072 28354
rect 414020 28290 414072 28296
rect 407120 24200 407172 24206
rect 407120 24142 407172 24148
rect 398840 22840 398892 22846
rect 398840 22782 398892 22788
rect 398852 2378 398880 22782
rect 407132 16574 407160 24142
rect 414032 16574 414060 28290
rect 416792 16574 416820 44814
rect 572720 43444 572772 43450
rect 572720 43386 572772 43392
rect 498200 42084 498252 42090
rect 498200 42026 498252 42032
rect 481640 40724 481692 40730
rect 481640 40666 481692 40672
rect 431960 37936 432012 37942
rect 431960 37878 432012 37884
rect 427820 17332 427872 17338
rect 427820 17274 427872 17280
rect 427832 16574 427860 17274
rect 431972 16574 432000 37878
rect 481652 16574 481680 40666
rect 498212 16574 498240 42026
rect 563060 39364 563112 39370
rect 563060 39306 563112 39312
rect 509240 28280 509292 28286
rect 509240 28222 509292 28228
rect 506480 17264 506532 17270
rect 506480 17206 506532 17212
rect 407132 16546 407252 16574
rect 414032 16546 414336 16574
rect 416792 16546 417464 16574
rect 427832 16546 428504 16574
rect 431972 16546 432092 16574
rect 481652 16546 481772 16574
rect 498212 16546 498976 16574
rect 403624 8152 403676 8158
rect 403624 8094 403676 8100
rect 398840 2372 398892 2378
rect 398840 2314 398892 2320
rect 400128 2372 400180 2378
rect 400128 2314 400180 2320
rect 400140 480 400168 2314
rect 403636 480 403664 8094
rect 407224 480 407252 16546
rect 410800 8084 410852 8090
rect 410800 8026 410852 8032
rect 410812 480 410840 8026
rect 414308 480 414336 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 420920 14544 420972 14550
rect 420920 14486 420972 14492
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 14486
rect 424968 8016 425020 8022
rect 424968 7958 425020 7964
rect 424980 480 425008 7958
rect 428476 480 428504 16546
rect 432064 480 432092 16546
rect 463976 15972 464028 15978
rect 463976 15914 464028 15920
rect 442632 13184 442684 13190
rect 442632 13126 442684 13132
rect 439136 7948 439188 7954
rect 439136 7890 439188 7896
rect 435548 3800 435600 3806
rect 435548 3742 435600 3748
rect 435560 480 435588 3742
rect 439148 480 439176 7890
rect 442644 480 442672 13126
rect 448520 10396 448572 10402
rect 448520 10338 448572 10344
rect 446220 7880 446272 7886
rect 446220 7822 446272 7828
rect 446232 480 446260 7822
rect 448532 3398 448560 10338
rect 453304 7812 453356 7818
rect 453304 7754 453356 7760
rect 448520 3392 448572 3398
rect 448520 3334 448572 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 453316 480 453344 7754
rect 460388 7744 460440 7750
rect 460388 7686 460440 7692
rect 456892 3732 456944 3738
rect 456892 3674 456944 3680
rect 456904 480 456932 3674
rect 460400 480 460428 7686
rect 463988 480 464016 15914
rect 478144 8968 478196 8974
rect 478144 8910 478196 8916
rect 467472 7676 467524 7682
rect 467472 7618 467524 7624
rect 467484 480 467512 7618
rect 474556 7608 474608 7614
rect 474556 7550 474608 7556
rect 471060 3664 471112 3670
rect 471060 3606 471112 3612
rect 471072 480 471100 3606
rect 474568 480 474596 7550
rect 478156 480 478184 8910
rect 481744 480 481772 16546
rect 495440 14476 495492 14482
rect 495440 14418 495492 14424
rect 492312 13116 492364 13122
rect 492312 13058 492364 13064
rect 488816 11756 488868 11762
rect 488816 11698 488868 11704
rect 484768 10328 484820 10334
rect 484768 10270 484820 10276
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 10270
rect 488828 480 488856 11698
rect 492324 480 492352 13058
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 354 495480 14418
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 502984 15904 503036 15910
rect 502984 15846 503036 15852
rect 502996 480 503024 15846
rect 506492 480 506520 17206
rect 509252 16574 509280 28222
rect 552020 24132 552072 24138
rect 552020 24074 552072 24080
rect 547880 18624 547932 18630
rect 547880 18566 547932 18572
rect 547892 16574 547920 18566
rect 552032 16574 552060 24074
rect 558920 22772 558972 22778
rect 558920 22714 558972 22720
rect 556160 21412 556212 21418
rect 556160 21354 556212 21360
rect 509252 16546 509648 16574
rect 547892 16546 548656 16574
rect 552032 16546 552704 16574
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 513564 5432 513616 5438
rect 513564 5374 513616 5380
rect 513576 480 513604 5374
rect 517152 5364 517204 5370
rect 517152 5306 517204 5312
rect 517164 480 517192 5306
rect 520740 5296 520792 5302
rect 520740 5238 520792 5244
rect 520752 480 520780 5238
rect 524236 5228 524288 5234
rect 524236 5170 524288 5176
rect 524248 480 524276 5170
rect 527824 5160 527876 5166
rect 527824 5102 527876 5108
rect 527836 480 527864 5102
rect 531320 5092 531372 5098
rect 531320 5034 531372 5040
rect 531332 480 531360 5034
rect 534908 5024 534960 5030
rect 534908 4966 534960 4972
rect 534920 480 534948 4966
rect 538404 4956 538456 4962
rect 538404 4898 538456 4904
rect 538416 480 538444 4898
rect 541992 4888 542044 4894
rect 541992 4830 542044 4836
rect 542004 480 542032 4830
rect 545488 4820 545540 4826
rect 545488 4762 545540 4768
rect 545500 480 545528 4762
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 552676 480 552704 16546
rect 556172 480 556200 21354
rect 558932 16574 558960 22714
rect 558932 16546 559328 16574
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 39306
rect 569960 26920 570012 26926
rect 569960 26862 570012 26868
rect 565820 25560 565872 25566
rect 565820 25502 565872 25508
rect 565832 16574 565860 25502
rect 569972 16574 570000 26862
rect 572732 16574 572760 43386
rect 576860 29640 576912 29646
rect 576860 29582 576912 29588
rect 576872 16574 576900 29582
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 565832 16546 566872 16574
rect 569972 16546 570368 16574
rect 572732 16546 573496 16574
rect 576872 16546 576992 16574
rect 566844 480 566872 16546
rect 570340 480 570368 16546
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 579986 7576 580042 7585
rect 579986 7511 580042 7520
rect 580000 6633 580028 7511
rect 579986 6624 580042 6633
rect 579986 6559 580042 6568
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 583404 480 583432 3470
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 2778 579964 2834 580000
rect 2778 579944 2780 579964
rect 2780 579944 2832 579964
rect 2832 579944 2834 579964
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527876 3478 527912
rect 3422 527856 3424 527876
rect 3424 527856 3476 527876
rect 3476 527856 3478 527876
rect 3422 514800 3478 514856
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 410488 3570 410544
rect 3422 306176 3478 306232
rect 3422 293120 3478 293176
rect 170862 685908 170918 685944
rect 170862 685888 170864 685908
rect 170864 685888 170916 685908
rect 170916 685888 170918 685908
rect 37830 636248 37886 636304
rect 36818 596808 36874 596864
rect 37002 596944 37058 597000
rect 38474 635296 38530 635352
rect 38014 632168 38070 632224
rect 37830 517384 37886 517440
rect 37738 516024 37794 516080
rect 37830 507864 37886 507920
rect 37738 488280 37794 488336
rect 38106 630672 38162 630728
rect 38014 513304 38070 513360
rect 38290 629312 38346 629368
rect 38198 627952 38254 628008
rect 38106 510992 38162 511048
rect 38290 509904 38346 509960
rect 38198 507864 38254 507920
rect 38566 610000 38622 610056
rect 38474 513984 38530 514040
rect 39854 597352 39910 597408
rect 38566 489912 38622 489968
rect 38474 479984 38530 480040
rect 39578 597080 39634 597136
rect 56414 597488 56470 597544
rect 63222 597488 63278 597544
rect 64234 597488 64290 597544
rect 64878 597488 64934 597544
rect 66810 597508 66866 597544
rect 66810 597488 66812 597508
rect 66812 597488 66864 597508
rect 66864 597488 66866 597508
rect 56414 597080 56470 597136
rect 56598 597080 56654 597136
rect 59358 597080 59414 597136
rect 67638 597488 67694 597544
rect 68926 597488 68982 597544
rect 69754 597488 69810 597544
rect 71686 597488 71742 597544
rect 73158 597488 73214 597544
rect 74446 597488 74502 597544
rect 74906 597488 74962 597544
rect 77206 597488 77262 597544
rect 78034 597488 78090 597544
rect 78586 597488 78642 597544
rect 81346 597488 81402 597544
rect 84198 597508 84254 597544
rect 84198 597488 84200 597508
rect 84200 597488 84252 597508
rect 84252 597488 84254 597508
rect 55402 596672 55458 596728
rect 68834 597352 68890 597408
rect 71318 597352 71374 597408
rect 71778 597352 71834 597408
rect 76010 597352 76066 597408
rect 77114 597352 77170 597408
rect 74446 570696 74502 570752
rect 71686 566344 71742 566400
rect 86866 597488 86922 597544
rect 88246 597488 88302 597544
rect 92478 597488 92534 597544
rect 93766 597488 93822 597544
rect 124126 597488 124182 597544
rect 129646 597488 129702 597544
rect 131026 597488 131082 597544
rect 133786 597488 133842 597544
rect 136546 597488 136602 597544
rect 142066 597488 142122 597544
rect 146206 597488 146262 597544
rect 82818 597352 82874 597408
rect 81438 597216 81494 597272
rect 85578 597216 85634 597272
rect 82818 596828 82874 596864
rect 82818 596808 82820 596828
rect 82820 596808 82872 596828
rect 82872 596808 82874 596828
rect 84106 596400 84162 596456
rect 86958 597216 87014 597272
rect 88338 597080 88394 597136
rect 89718 597080 89774 597136
rect 91190 596536 91246 596592
rect 91098 596420 91154 596456
rect 91098 596400 91100 596420
rect 91100 596400 91152 596420
rect 91152 596400 91154 596420
rect 91006 596264 91062 596320
rect 108946 597352 109002 597408
rect 117226 597352 117282 597408
rect 121366 597352 121422 597408
rect 95238 597236 95294 597272
rect 95238 597216 95240 597236
rect 95240 597216 95292 597236
rect 95292 597216 95294 597236
rect 96618 597100 96674 597136
rect 96618 597080 96620 597100
rect 96620 597080 96672 597100
rect 96672 597080 96674 597100
rect 102046 596672 102102 596728
rect 94042 596536 94098 596592
rect 96526 596400 96582 596456
rect 99286 596400 99342 596456
rect 106186 596536 106242 596592
rect 114466 597216 114522 597272
rect 111706 596944 111762 597000
rect 118606 596964 118662 597000
rect 118606 596944 118608 596964
rect 118608 596944 118660 596964
rect 118660 596944 118662 596964
rect 126886 597080 126942 597136
rect 139306 597100 139362 597136
rect 139306 597080 139308 597100
rect 139308 597080 139360 597100
rect 139360 597080 139362 597100
rect 170862 565800 170918 565856
rect 146206 565392 146262 565448
rect 129646 565256 129702 565312
rect 93766 565120 93822 565176
rect 68926 564984 68982 565040
rect 56046 479576 56102 479632
rect 72330 478644 72386 478680
rect 72330 478624 72332 478644
rect 72332 478624 72384 478644
rect 72384 478624 72386 478644
rect 74630 478624 74686 478680
rect 73158 478508 73214 478544
rect 73158 478488 73160 478508
rect 73160 478488 73212 478508
rect 73212 478488 73214 478508
rect 63222 477400 63278 477456
rect 64234 477400 64290 477456
rect 64878 477400 64934 477456
rect 66534 477400 66590 477456
rect 67638 477400 67694 477456
rect 68742 477400 68798 477456
rect 70214 477420 70270 477456
rect 70214 477400 70216 477420
rect 70216 477400 70268 477420
rect 70268 477400 70270 477420
rect 59450 477264 59506 477320
rect 60738 477264 60794 477320
rect 58162 476856 58218 476912
rect 70858 477436 70860 477456
rect 70860 477436 70912 477456
rect 70912 477436 70914 477456
rect 70858 477400 70914 477436
rect 57886 476740 57942 476776
rect 57886 476720 57888 476740
rect 57888 476720 57940 476740
rect 57940 476720 57942 476740
rect 76930 478488 76986 478544
rect 75826 478372 75882 478408
rect 75826 478352 75828 478372
rect 75828 478352 75880 478372
rect 75880 478352 75882 478372
rect 78126 477400 78182 477456
rect 79506 478236 79562 478272
rect 79506 478216 79508 478236
rect 79508 478216 79560 478236
rect 79560 478216 79562 478236
rect 80610 478116 80612 478136
rect 80612 478116 80664 478136
rect 80664 478116 80666 478136
rect 80610 478080 80666 478116
rect 81346 477400 81402 477456
rect 81806 477400 81862 477456
rect 68926 476176 68982 476232
rect 71686 476176 71742 476232
rect 74446 476176 74502 476232
rect 77206 476176 77262 476232
rect 78586 476176 78642 476232
rect 86314 477536 86370 477592
rect 82818 477400 82874 477456
rect 84106 477400 84162 477456
rect 85302 477400 85358 477456
rect 82726 476176 82782 476232
rect 84014 476584 84070 476640
rect 86866 477400 86922 477456
rect 87602 477436 87604 477456
rect 87604 477436 87656 477456
rect 87656 477436 87658 477456
rect 87602 477400 87658 477436
rect 88246 477400 88302 477456
rect 88706 477400 88762 477456
rect 89718 477400 89774 477456
rect 91190 477400 91246 477456
rect 92202 477400 92258 477456
rect 93030 477400 93086 477456
rect 94410 477400 94466 477456
rect 95790 477400 95846 477456
rect 96986 477400 97042 477456
rect 91006 476448 91062 476504
rect 93766 476448 93822 476504
rect 95974 476448 96030 476504
rect 95974 476176 96030 476232
rect 96526 476176 96582 476232
rect 99286 476176 99342 476232
rect 102046 476176 102102 476232
rect 104806 476176 104862 476232
rect 106186 476176 106242 476232
rect 108946 476176 109002 476232
rect 111706 476176 111762 476232
rect 114466 476176 114522 476232
rect 117226 476176 117282 476232
rect 118606 476176 118662 476232
rect 121366 476176 121422 476232
rect 124126 476176 124182 476232
rect 126886 476176 126942 476232
rect 129646 476176 129702 476232
rect 131026 476176 131082 476232
rect 133786 476176 133842 476232
rect 136546 476176 136602 476232
rect 139306 476176 139362 476232
rect 142066 476176 142122 476232
rect 143446 476176 143502 476232
rect 146206 476176 146262 476232
rect 111706 445168 111762 445224
rect 108946 445032 109002 445088
rect 93766 444896 93822 444952
rect 170862 445712 170918 445768
rect 74446 443536 74502 443592
rect 38474 397296 38530 397352
rect 38474 395392 38530 395448
rect 37738 368328 37794 368384
rect 38198 368328 38254 368384
rect 38382 367512 38438 367568
rect 39026 393488 39082 393544
rect 38842 392264 38898 392320
rect 38750 389408 38806 389464
rect 38658 387776 38714 387832
rect 38566 369824 38622 369880
rect 38934 390632 38990 390688
rect 61382 358128 61438 358184
rect 64326 358128 64382 358184
rect 56506 357312 56562 357368
rect 59266 357312 59322 357368
rect 60646 357312 60702 357368
rect 58622 357176 58678 357232
rect 62026 357312 62082 357368
rect 63406 357312 63462 357368
rect 67546 357312 67602 357368
rect 68834 357312 68890 357368
rect 70306 357312 70362 357368
rect 71686 357312 71742 357368
rect 73066 357312 73122 357368
rect 74354 357312 74410 357368
rect 75826 357312 75882 357368
rect 76010 357312 76066 357368
rect 78586 357312 78642 357368
rect 79966 357312 80022 357368
rect 81346 357312 81402 357368
rect 86866 357312 86922 357368
rect 88246 357312 88302 357368
rect 91006 357312 91062 357368
rect 93398 357312 93454 357368
rect 96526 357312 96582 357368
rect 99286 357312 99342 357368
rect 102046 357312 102102 357368
rect 106186 357312 106242 357368
rect 66166 356088 66222 356144
rect 68926 357040 68982 357096
rect 68926 356108 68982 356144
rect 68926 356088 68928 356108
rect 68928 356088 68980 356108
rect 68980 356088 68982 356108
rect 71594 357176 71650 357232
rect 74078 357176 74134 357232
rect 77022 357176 77078 357232
rect 78494 357176 78550 357232
rect 77206 356360 77262 356416
rect 81254 357176 81310 357232
rect 84106 356632 84162 356688
rect 104806 356088 104862 356144
rect 144642 355272 144698 355328
rect 138754 353912 138810 353968
rect 3330 267144 3386 267200
rect 2962 254088 3018 254144
rect 3330 241032 3386 241088
rect 3054 214920 3110 214976
rect 3330 188808 3386 188864
rect 3054 162832 3110 162888
rect 3330 149776 3386 149832
rect 3330 136720 3386 136776
rect 3330 110608 3386 110664
rect 3330 97552 3386 97608
rect 3790 201864 3846 201920
rect 3698 84632 3754 84688
rect 3606 71576 3662 71632
rect 3514 58520 3570 58576
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 32408 3478 32464
rect 3422 19352 3478 19408
rect 125506 281696 125562 281752
rect 126886 281832 126942 281888
rect 127760 280200 127816 280256
rect 128726 281560 128782 281616
rect 133970 290400 134026 290456
rect 136454 284824 136510 284880
rect 142802 352552 142858 352608
rect 141330 351056 141386 351112
rect 140594 349696 140650 349752
rect 140962 290536 141018 290592
rect 143906 337320 143962 337376
rect 145010 342896 145066 342952
rect 145746 327664 145802 327720
rect 148598 282104 148654 282160
rect 175186 281832 175242 281888
rect 175186 280744 175242 280800
rect 175922 281696 175978 281752
rect 175922 280880 175978 280936
rect 177210 596944 177266 597000
rect 177486 290808 177542 290864
rect 177670 290672 177726 290728
rect 178130 282784 178186 282840
rect 178498 679088 178554 679144
rect 178498 560224 178554 560280
rect 178498 439184 178554 439240
rect 179050 560224 179106 560280
rect 179050 559136 179106 559192
rect 180154 487192 180210 487248
rect 181810 287272 181866 287328
rect 178774 281696 178830 281752
rect 183466 282104 183522 282160
rect 185582 281560 185638 281616
rect 186226 281560 186282 281616
rect 187698 287136 187754 287192
rect 189906 287408 189962 287464
rect 188986 281968 189042 282024
rect 191286 281832 191342 281888
rect 235170 700712 235226 700768
rect 267646 700576 267702 700632
rect 300122 700440 300178 700496
rect 332506 700304 332562 700360
rect 350998 685908 351054 685944
rect 350998 685888 351000 685908
rect 351000 685888 351052 685908
rect 351052 685888 351054 685908
rect 358818 678952 358874 679008
rect 217230 636792 217286 636848
rect 217138 635840 217194 635896
rect 216678 608232 216734 608288
rect 213550 597352 213606 597408
rect 211066 596944 211122 597000
rect 210698 477400 210754 477456
rect 210422 477264 210478 477320
rect 203614 290944 203670 291000
rect 210422 476584 210478 476640
rect 208674 294480 208730 294536
rect 209226 282784 209282 282840
rect 210514 476448 210570 476504
rect 210882 477128 210938 477184
rect 210698 476312 210754 476368
rect 210698 282784 210754 282840
rect 213366 477264 213422 477320
rect 213274 476992 213330 477048
rect 213182 476856 213238 476912
rect 212354 359488 212410 359544
rect 211526 282784 211582 282840
rect 211618 282648 211674 282704
rect 213366 476720 213422 476776
rect 213274 355952 213330 356008
rect 213642 594496 213698 594552
rect 213550 358264 213606 358320
rect 213734 594360 213790 594416
rect 213642 355816 213698 355872
rect 213826 594224 213882 594280
rect 213734 355680 213790 355736
rect 213918 567180 213974 567216
rect 213918 567160 213920 567180
rect 213920 567160 213972 567180
rect 213972 567160 213974 567180
rect 214470 476448 214526 476504
rect 216586 596672 216642 596728
rect 214654 476312 214710 476368
rect 213826 355544 213882 355600
rect 213090 293120 213146 293176
rect 213642 282648 213698 282704
rect 214286 285232 214342 285288
rect 214470 285096 214526 285152
rect 214746 285368 214802 285424
rect 216126 474000 216182 474056
rect 216770 516160 216826 516216
rect 217874 633664 217930 633720
rect 217690 632712 217746 632768
rect 217598 630944 217654 631000
rect 217506 629856 217562 629912
rect 217414 628088 217470 628144
rect 217230 516840 217286 516896
rect 217230 516160 217286 516216
rect 216954 515888 217010 515944
rect 217138 515888 217194 515944
rect 217046 513712 217102 513768
rect 217138 512760 217194 512816
rect 217046 479984 217102 480040
rect 217046 478896 217102 478952
rect 216954 391856 217010 391912
rect 216954 391040 217010 391096
rect 216862 390496 216918 390552
rect 216678 369960 216734 370016
rect 216862 369824 216918 369880
rect 216862 368328 216918 368384
rect 216586 358536 216642 358592
rect 215022 284960 215078 285016
rect 215850 282784 215906 282840
rect 216218 282784 216274 282840
rect 217138 392808 217194 392864
rect 217782 610000 217838 610056
rect 217690 512760 217746 512816
rect 217598 510992 217654 511048
rect 217506 509904 217562 509960
rect 217414 508136 217470 508192
rect 258078 599528 258134 599584
rect 277306 599528 277362 599584
rect 235998 597488 236054 597544
rect 236182 597488 236238 597544
rect 237378 597488 237434 597544
rect 243082 597488 243138 597544
rect 244278 597488 244334 597544
rect 245474 597488 245530 597544
rect 246486 597488 246542 597544
rect 247038 597488 247094 597544
rect 248418 597488 248474 597544
rect 249798 597488 249854 597544
rect 252098 597488 252154 597544
rect 253478 597488 253534 597544
rect 254582 597488 254638 597544
rect 255410 597488 255466 597544
rect 256698 597488 256754 597544
rect 219990 597080 220046 597136
rect 217874 513712 217930 513768
rect 217782 489912 217838 489968
rect 218426 488008 218482 488064
rect 217506 477128 217562 477184
rect 217966 477128 218022 477184
rect 217506 476584 217562 476640
rect 217322 395936 217378 395992
rect 217230 391856 217286 391912
rect 217230 388184 217286 388240
rect 217690 396888 217746 396944
rect 217414 388184 217470 388240
rect 217414 368056 217470 368112
rect 217874 390496 217930 390552
rect 217874 389952 217930 390008
rect 218150 474680 218206 474736
rect 218150 393896 218206 393952
rect 218886 477264 218942 477320
rect 218978 476992 219034 477048
rect 219070 476856 219126 476912
rect 219254 477400 219310 477456
rect 218886 474136 218942 474192
rect 218610 393760 218666 393816
rect 218518 392808 218574 392864
rect 218518 368328 218574 368384
rect 218794 395936 218850 395992
rect 217690 282784 217746 282840
rect 218426 282784 218482 282840
rect 219346 358400 219402 358456
rect 219898 474680 219954 474736
rect 238758 596828 238814 596864
rect 238758 596808 238760 596828
rect 238760 596808 238812 596828
rect 238812 596808 238814 596828
rect 240138 596808 240194 596864
rect 241518 596808 241574 596864
rect 247130 596808 247186 596864
rect 247038 566480 247094 566536
rect 249890 596808 249946 596864
rect 252190 596808 252246 596864
rect 260838 597488 260894 597544
rect 263598 597488 263654 597544
rect 264978 597488 265034 597544
rect 267738 597488 267794 597544
rect 270498 597488 270554 597544
rect 276018 597488 276074 597544
rect 262218 597352 262274 597408
rect 259550 596672 259606 596728
rect 259458 596536 259514 596592
rect 263690 597352 263746 597408
rect 263598 594496 263654 594552
rect 266358 597352 266414 597408
rect 265070 596828 265126 596864
rect 265070 596808 265072 596828
rect 265072 596808 265124 596828
rect 265124 596808 265126 596828
rect 266358 596436 266360 596456
rect 266360 596436 266412 596456
rect 266412 596436 266414 596456
rect 266358 596400 266414 596436
rect 264978 594360 265034 594416
rect 270406 597352 270462 597408
rect 270406 597080 270462 597136
rect 267922 596672 267978 596728
rect 269118 596692 269174 596728
rect 269118 596672 269120 596692
rect 269120 596672 269172 596692
rect 269172 596672 269174 596692
rect 267738 594224 267794 594280
rect 274638 597236 274694 597272
rect 274638 597216 274640 597236
rect 274640 597216 274692 597236
rect 274692 597216 274694 597236
rect 270590 597080 270646 597136
rect 273258 597080 273314 597136
rect 280158 597488 280214 597544
rect 282918 597488 282974 597544
rect 285678 597488 285734 597544
rect 289818 597488 289874 597544
rect 292578 597488 292634 597544
rect 277306 596944 277362 597000
rect 271878 596420 271934 596456
rect 271878 596400 271880 596420
rect 271880 596400 271932 596420
rect 271932 596400 271934 596420
rect 273258 596264 273314 596320
rect 270498 594088 270554 594144
rect 287058 597080 287114 597136
rect 326986 596944 327042 597000
rect 311806 596808 311862 596864
rect 321466 596808 321522 596864
rect 324226 596828 324282 596864
rect 324226 596808 324228 596828
rect 324228 596808 324280 596828
rect 324280 596808 324282 596828
rect 356794 596808 356850 596864
rect 314566 596672 314622 596728
rect 318706 596692 318762 596728
rect 318706 596672 318708 596692
rect 318708 596672 318760 596692
rect 318760 596672 318762 596692
rect 315946 596556 316002 596592
rect 315946 596536 315948 596556
rect 315948 596536 316000 596556
rect 316000 596536 316002 596556
rect 306102 596400 306158 596456
rect 309046 596420 309102 596456
rect 309046 596400 309048 596420
rect 309048 596400 309100 596420
rect 309100 596400 309102 596420
rect 296350 596264 296406 596320
rect 303526 596284 303582 596320
rect 303526 596264 303528 596284
rect 303528 596264 303580 596284
rect 303580 596264 303582 596284
rect 282918 593952 282974 594008
rect 351090 565800 351146 565856
rect 235998 479576 236054 479632
rect 243174 477400 243230 477456
rect 244278 477400 244334 477456
rect 245474 477400 245530 477456
rect 245934 477400 245990 477456
rect 247130 477400 247186 477456
rect 248602 477400 248658 477456
rect 250074 477400 250130 477456
rect 251270 477400 251326 477456
rect 252374 477436 252376 477456
rect 252376 477436 252428 477456
rect 252428 477436 252430 477456
rect 252374 477400 252430 477436
rect 253386 477400 253442 477456
rect 254490 477400 254546 477456
rect 255318 477420 255374 477456
rect 255318 477400 255320 477420
rect 255320 477400 255372 477420
rect 255372 477400 255374 477420
rect 256974 477400 257030 477456
rect 260838 477420 260894 477456
rect 260838 477400 260840 477420
rect 260840 477400 260892 477420
rect 260892 477400 260894 477420
rect 266358 477400 266414 477456
rect 269118 477436 269120 477456
rect 269120 477436 269172 477456
rect 269172 477436 269174 477456
rect 269118 477400 269174 477436
rect 278778 477420 278834 477456
rect 278778 477400 278780 477420
rect 278780 477400 278832 477420
rect 278832 477400 278834 477420
rect 259366 477264 259422 477320
rect 260838 477264 260894 477320
rect 263598 477284 263654 477320
rect 263598 477264 263600 477284
rect 263600 477264 263652 477284
rect 263652 477264 263654 477284
rect 255318 476856 255374 476912
rect 247038 476176 247094 476232
rect 249798 476176 249854 476232
rect 252558 476176 252614 476232
rect 258262 476176 258318 476232
rect 271878 477264 271934 477320
rect 276018 477264 276074 477320
rect 277674 477284 277730 477320
rect 277674 477264 277676 477284
rect 277676 477264 277728 477284
rect 277728 477264 277730 477284
rect 262218 476856 262274 476912
rect 264978 476992 265034 477048
rect 270498 477012 270554 477048
rect 270498 476992 270500 477012
rect 270500 476992 270552 477012
rect 270552 476992 270554 477012
rect 270498 476856 270554 476912
rect 273258 477148 273314 477184
rect 273258 477128 273260 477148
rect 273260 477128 273312 477148
rect 273312 477128 273314 477148
rect 274638 477128 274694 477184
rect 311806 477128 311862 477184
rect 277582 476992 277638 477048
rect 285678 476992 285734 477048
rect 266358 476720 266414 476776
rect 263690 476584 263746 476640
rect 268198 476604 268254 476640
rect 268198 476584 268200 476604
rect 268200 476584 268252 476604
rect 268252 476584 268254 476604
rect 255318 474136 255374 474192
rect 260838 476176 260894 476232
rect 263598 476176 263654 476232
rect 264978 476176 265034 476232
rect 268014 476176 268070 476232
rect 258262 474000 258318 474056
rect 273258 476856 273314 476912
rect 273258 476176 273314 476232
rect 276018 476176 276074 476232
rect 280158 476176 280214 476232
rect 282918 476176 282974 476232
rect 287702 476720 287758 476776
rect 302146 476720 302202 476776
rect 289818 476448 289874 476504
rect 299386 476312 299442 476368
rect 292578 476176 292634 476232
rect 296258 476176 296314 476232
rect 309046 476584 309102 476640
rect 306102 476448 306158 476504
rect 324226 476992 324282 477048
rect 326986 476992 327042 477048
rect 321466 476856 321522 476912
rect 315946 476720 316002 476776
rect 318706 476740 318762 476776
rect 318706 476720 318708 476740
rect 318708 476720 318760 476740
rect 318760 476720 318762 476740
rect 314566 476604 314622 476640
rect 314566 476584 314568 476604
rect 314568 476584 314620 476604
rect 314620 476584 314622 476604
rect 303526 476332 303582 476368
rect 303526 476312 303528 476332
rect 303528 476312 303580 476332
rect 303580 476312 303582 476332
rect 351090 445712 351146 445768
rect 221922 359896 221978 359952
rect 219990 357992 220046 358048
rect 220082 311072 220138 311128
rect 220266 282784 220322 282840
rect 223762 358672 223818 358728
rect 228178 358536 228234 358592
rect 224222 358400 224278 358456
rect 225234 356632 225290 356688
rect 227074 290944 227130 291000
rect 263874 359624 263930 359680
rect 253202 359488 253258 359544
rect 253202 359216 253258 359272
rect 235998 358556 236054 358592
rect 235998 358536 236000 358556
rect 236000 358536 236052 358556
rect 236052 358536 236054 358556
rect 234066 358400 234122 358456
rect 232226 358264 232282 358320
rect 229282 298696 229338 298752
rect 233330 297336 233386 297392
rect 234434 324944 234490 325000
rect 238022 357176 238078 357232
rect 237010 356224 237066 356280
rect 236274 355816 236330 355872
rect 237010 351192 237066 351248
rect 237378 348336 237434 348392
rect 238758 357040 238814 357096
rect 238482 304136 238538 304192
rect 243542 357312 243598 357368
rect 240230 355952 240286 356008
rect 240322 355680 240378 355736
rect 244922 356904 244978 356960
rect 245106 356904 245162 356960
rect 244002 355544 244058 355600
rect 245566 356632 245622 356688
rect 246854 356360 246910 356416
rect 245106 356088 245162 356144
rect 247222 357312 247278 357368
rect 248694 357312 248750 357368
rect 249982 357312 250038 357368
rect 247130 356496 247186 356552
rect 247314 355408 247370 355464
rect 250074 356632 250130 356688
rect 249522 293528 249578 293584
rect 248970 282512 249026 282568
rect 250626 358128 250682 358184
rect 251270 357312 251326 357368
rect 252650 357312 252706 357368
rect 251362 354048 251418 354104
rect 252282 356632 252338 356688
rect 253386 356496 253442 356552
rect 252834 290808 252890 290864
rect 253938 357992 253994 358048
rect 254582 357312 254638 357368
rect 255410 357312 255466 357368
rect 255042 351328 255098 351384
rect 255778 356632 255834 356688
rect 256146 290672 256202 290728
rect 255594 285368 255650 285424
rect 257342 357312 257398 357368
rect 258170 357312 258226 357368
rect 257986 354184 258042 354240
rect 258814 356632 258870 356688
rect 258906 285232 258962 285288
rect 260562 359216 260618 359272
rect 260194 356632 260250 356688
rect 260102 356360 260158 356416
rect 260838 357312 260894 357368
rect 262126 357348 262128 357368
rect 262128 357348 262180 357368
rect 262180 357348 262182 357368
rect 262126 357312 262182 357348
rect 262770 357332 262826 357368
rect 262770 357312 262772 357332
rect 262772 357312 262824 357332
rect 262824 357312 262826 357332
rect 262770 289040 262826 289096
rect 262218 285096 262274 285152
rect 263690 357312 263746 357368
rect 263966 357312 264022 357368
rect 266634 359352 266690 359408
rect 265714 357312 265770 357368
rect 266450 357312 266506 357368
rect 264978 356496 265034 356552
rect 265530 284960 265586 285016
rect 267554 357312 267610 357368
rect 267738 357312 267794 357368
rect 268566 357312 268622 357368
rect 269762 357312 269818 357368
rect 267922 354320 267978 354376
rect 269026 287816 269082 287872
rect 270590 357312 270646 357368
rect 271142 357312 271198 357368
rect 272154 357312 272210 357368
rect 271970 287680 272026 287736
rect 273350 357312 273406 357368
rect 273350 356088 273406 356144
rect 276018 358128 276074 358184
rect 274546 357312 274602 357368
rect 275926 357312 275982 357368
rect 274178 354456 274234 354512
rect 277030 357312 277086 357368
rect 277398 356088 277454 356144
rect 285218 359488 285274 359544
rect 282274 359352 282330 359408
rect 280158 356088 280214 356144
rect 282918 357312 282974 357368
rect 285678 357312 285734 357368
rect 287058 357312 287114 357368
rect 289910 357312 289966 357368
rect 292578 357312 292634 357368
rect 292946 293392 293002 293448
rect 294050 357992 294106 358048
rect 295338 357312 295394 357368
rect 296994 357856 297050 357912
rect 298190 357312 298246 357368
rect 299938 358264 299994 358320
rect 308770 358536 308826 358592
rect 300858 358128 300914 358184
rect 301042 358128 301098 358184
rect 301042 357856 301098 357912
rect 302238 357312 302294 357368
rect 304998 357312 305054 357368
rect 305826 358400 305882 358456
rect 307758 357312 307814 357368
rect 310518 357312 310574 357368
rect 313278 357312 313334 357368
rect 313554 293256 313610 293312
rect 325698 358672 325754 358728
rect 314750 357312 314806 357368
rect 317418 357312 317474 357368
rect 320178 357312 320234 357368
rect 316682 342896 316738 342952
rect 322938 356088 322994 356144
rect 356702 476720 356758 476776
rect 356610 357992 356666 358048
rect 356886 476992 356942 477048
rect 357070 476856 357126 476912
rect 357530 358264 357586 358320
rect 358818 560224 358874 560280
rect 357714 358400 357770 358456
rect 357622 358128 357678 358184
rect 358818 439184 358874 439240
rect 315762 282240 315818 282296
rect 123850 279520 123906 279576
rect 123712 279248 123768 279304
rect 318246 271904 318302 271960
rect 318154 233824 318210 233880
rect 319626 287408 319682 287464
rect 320822 287272 320878 287328
rect 319810 282104 319866 282160
rect 318062 232464 318118 232520
rect 318062 230560 318118 230616
rect 318154 229064 318210 229120
rect 3422 6432 3478 6488
rect 359094 358536 359150 358592
rect 359738 560224 359794 560280
rect 359738 559136 359794 559192
rect 389822 597216 389878 597272
rect 370502 477128 370558 477184
rect 389730 593952 389786 594008
rect 390098 594360 390154 594416
rect 390466 594224 390522 594280
rect 390282 594088 390338 594144
rect 494794 700440 494850 700496
rect 527178 700304 527234 700360
rect 397458 699760 397514 699816
rect 530950 685908 531006 685944
rect 530950 685888 530952 685908
rect 530952 685888 531004 685908
rect 531004 685888 531006 685908
rect 397274 636792 397330 636848
rect 396906 635840 396962 635896
rect 396630 632712 396686 632768
rect 392674 597352 392730 597408
rect 392858 596400 392914 596456
rect 392674 351328 392730 351384
rect 393962 356632 394018 356688
rect 394514 356632 394570 356688
rect 393870 356496 393926 356552
rect 394514 356360 394570 356416
rect 396446 516160 396502 516216
rect 396538 514800 396594 514856
rect 396814 628088 396870 628144
rect 396722 610000 396778 610056
rect 396630 512760 396686 512816
rect 396998 633664 397054 633720
rect 396906 515888 396962 515944
rect 396906 514800 396962 514856
rect 397090 630944 397146 631000
rect 396998 513712 397054 513768
rect 396998 512760 397054 512816
rect 396906 510448 396962 510504
rect 396906 509904 396962 509960
rect 396814 508136 396870 508192
rect 396722 489912 396778 489968
rect 396630 396888 396686 396944
rect 396538 395936 396594 395992
rect 396630 394576 396686 394632
rect 396630 393760 396686 393816
rect 396446 369960 396502 370016
rect 396538 368056 396594 368112
rect 397182 608232 397238 608288
rect 397090 510992 397146 511048
rect 396998 392808 397054 392864
rect 396906 389952 396962 390008
rect 396814 388184 396870 388240
rect 396722 369960 396778 370016
rect 396722 368328 396778 368384
rect 397366 629856 397422 629912
rect 397274 516840 397330 516896
rect 397274 516160 397330 516216
rect 435914 599528 435970 599584
rect 415398 597488 415454 597544
rect 416778 597488 416834 597544
rect 418158 597488 418214 597544
rect 419538 597488 419594 597544
rect 420918 597488 420974 597544
rect 423126 597488 423182 597544
rect 424966 597488 425022 597544
rect 425610 597488 425666 597544
rect 426530 597488 426586 597544
rect 427634 597488 427690 597544
rect 428002 597488 428058 597544
rect 429198 597488 429254 597544
rect 430578 597488 430634 597544
rect 433338 597488 433394 597544
rect 434534 597488 434590 597544
rect 397366 510448 397422 510504
rect 397182 488280 397238 488336
rect 397182 487328 397238 487384
rect 397090 391040 397146 391096
rect 398562 477264 398618 477320
rect 398102 476584 398158 476640
rect 397826 474272 397882 474328
rect 398010 474000 398066 474056
rect 397182 356768 397238 356824
rect 397918 354320 397974 354376
rect 398286 476312 398342 476368
rect 398194 474408 398250 474464
rect 398470 474136 398526 474192
rect 398930 357312 398986 357368
rect 399390 357176 399446 357232
rect 398930 356224 398986 356280
rect 398470 354456 398526 354512
rect 398286 354184 398342 354240
rect 398102 354048 398158 354104
rect 419538 596672 419594 596728
rect 427818 596672 427874 596728
rect 427818 571920 427874 571976
rect 430670 596672 430726 596728
rect 431958 596672 432014 596728
rect 430578 570560 430634 570616
rect 434718 597488 434774 597544
rect 451094 599392 451150 599448
rect 437110 597488 437166 597544
rect 437478 597488 437534 597544
rect 438858 597488 438914 597544
rect 441986 597488 442042 597544
rect 442998 597488 443054 597544
rect 443642 597488 443698 597544
rect 444378 597488 444434 597544
rect 445758 597488 445814 597544
rect 447138 597488 447194 597544
rect 449898 597488 449954 597544
rect 433430 596672 433486 596728
rect 440330 597080 440386 597136
rect 438858 596672 438914 596728
rect 441618 596944 441674 597000
rect 442998 594496 443054 594552
rect 445850 596944 445906 597000
rect 447230 596944 447286 597000
rect 448518 596944 448574 597000
rect 448518 596284 448574 596320
rect 448518 596264 448520 596284
rect 448520 596264 448572 596284
rect 448572 596264 448574 596284
rect 462318 597488 462374 597544
rect 465078 597488 465134 597544
rect 467838 597488 467894 597544
rect 473358 597488 473414 597544
rect 474738 597488 474794 597544
rect 477498 597488 477554 597544
rect 483018 597488 483074 597544
rect 485778 597488 485834 597544
rect 488538 597488 488594 597544
rect 495438 597488 495494 597544
rect 498198 597488 498254 597544
rect 500958 597488 501014 597544
rect 452658 597352 452714 597408
rect 454038 596964 454094 597000
rect 454038 596944 454040 596964
rect 454040 596944 454092 596964
rect 454092 596944 454094 596964
rect 455418 596944 455474 597000
rect 449990 596420 450046 596456
rect 449990 596400 449992 596420
rect 449992 596400 450044 596420
rect 450044 596400 450046 596420
rect 451094 596400 451150 596456
rect 451278 596400 451334 596456
rect 456798 596264 456854 596320
rect 462318 594360 462374 594416
rect 465078 594224 465134 594280
rect 470598 596264 470654 596320
rect 467838 594088 467894 594144
rect 470598 593952 470654 594008
rect 480258 596944 480314 597000
rect 492678 596672 492734 596728
rect 489918 596264 489974 596320
rect 502338 596944 502394 597000
rect 505098 596808 505154 596864
rect 505098 592592 505154 592648
rect 538218 678952 538274 679008
rect 530950 565836 530952 565856
rect 530952 565836 531004 565856
rect 531004 565836 531006 565856
rect 530950 565800 531006 565836
rect 433338 563624 433394 563680
rect 415398 477400 415454 477456
rect 416778 477400 416834 477456
rect 418158 477400 418214 477456
rect 419538 477400 419594 477456
rect 420918 477400 420974 477456
rect 423126 477400 423182 477456
rect 424138 477400 424194 477456
rect 425518 477400 425574 477456
rect 419538 476448 419594 476504
rect 426622 477400 426678 477456
rect 427726 477400 427782 477456
rect 428554 478352 428610 478408
rect 430118 478372 430174 478408
rect 430118 478352 430120 478372
rect 430120 478352 430172 478372
rect 430172 478352 430174 478372
rect 431314 478236 431370 478272
rect 431314 478216 431316 478236
rect 431316 478216 431368 478236
rect 431368 478216 431370 478236
rect 432510 478216 432566 478272
rect 433430 477436 433432 477456
rect 433432 477436 433484 477456
rect 433484 477436 433486 477456
rect 433430 477400 433486 477436
rect 434534 477436 434536 477456
rect 434536 477436 434588 477456
rect 434588 477436 434590 477456
rect 434534 477400 434590 477436
rect 433338 476448 433394 476504
rect 427818 476176 427874 476232
rect 430578 476176 430634 476232
rect 399574 357040 399630 357096
rect 435730 477400 435786 477456
rect 436834 477400 436890 477456
rect 438122 477400 438178 477456
rect 442998 477400 443054 477456
rect 447138 477400 447194 477456
rect 448518 477420 448574 477456
rect 448518 477400 448520 477420
rect 448520 477400 448572 477420
rect 448572 477400 448574 477420
rect 438858 477128 438914 477184
rect 440238 476992 440294 477048
rect 441618 476856 441674 476912
rect 452658 477400 452714 477456
rect 444194 477128 444250 477184
rect 444378 477128 444434 477184
rect 445758 477148 445814 477184
rect 445758 477128 445760 477148
rect 445760 477128 445812 477148
rect 445812 477128 445814 477148
rect 448518 477164 448520 477184
rect 448520 477164 448572 477184
rect 448572 477164 448574 477184
rect 448518 477128 448574 477164
rect 451370 477128 451426 477184
rect 458178 477128 458234 477184
rect 462318 477128 462374 477184
rect 445666 477028 445668 477048
rect 445668 477028 445720 477048
rect 445720 477028 445722 477048
rect 445666 476992 445722 477028
rect 446402 476992 446458 477048
rect 454038 477012 454094 477048
rect 454038 476992 454040 477012
rect 454040 476992 454092 477012
rect 454092 476992 454094 477012
rect 456798 476992 456854 477048
rect 455418 476876 455474 476912
rect 455418 476856 455420 476876
rect 455420 476856 455472 476876
rect 455472 476856 455474 476876
rect 456890 476856 456946 476912
rect 446402 476584 446458 476640
rect 441986 476468 442042 476504
rect 441986 476448 441988 476468
rect 441988 476448 442040 476468
rect 442040 476448 442042 476468
rect 442998 476448 443054 476504
rect 449898 476448 449954 476504
rect 445758 476176 445814 476232
rect 447138 476176 447194 476232
rect 449898 476176 449954 476232
rect 442998 474544 443054 474600
rect 483018 476856 483074 476912
rect 474738 476448 474794 476504
rect 477498 476448 477554 476504
rect 465078 476176 465134 476232
rect 467838 476176 467894 476232
rect 470782 476176 470838 476232
rect 473358 476176 473414 476232
rect 462318 474408 462374 474464
rect 467838 474272 467894 474328
rect 470782 474136 470838 474192
rect 473358 474000 473414 474056
rect 480534 476176 480590 476232
rect 490470 476720 490526 476776
rect 498198 476720 498254 476776
rect 485778 476176 485834 476232
rect 488538 476176 488594 476232
rect 492678 476176 492734 476232
rect 495438 476176 495494 476232
rect 502338 476312 502394 476368
rect 500958 476176 501014 476232
rect 505098 476176 505154 476232
rect 430578 461488 430634 461544
rect 427818 460128 427874 460184
rect 530490 446392 530546 446448
rect 400126 444216 400182 444272
rect 416042 358128 416098 358184
rect 488538 358128 488594 358184
rect 423126 357348 423128 357368
rect 423128 357348 423180 357368
rect 423180 357348 423182 357368
rect 423126 357312 423182 357348
rect 399666 356904 399722 356960
rect 424966 357312 425022 357368
rect 425426 357312 425482 357368
rect 426898 357312 426954 357368
rect 427634 357312 427690 357368
rect 427818 357312 427874 357368
rect 428554 357312 428610 357368
rect 430026 357312 430082 357368
rect 430578 357312 430634 357368
rect 431958 357312 432014 357368
rect 433338 357312 433394 357368
rect 430670 357176 430726 357232
rect 434718 357312 434774 357368
rect 436834 357312 436890 357368
rect 437478 357312 437534 357368
rect 440238 357312 440294 357368
rect 444286 357312 444342 357368
rect 445850 357312 445906 357368
rect 447230 357312 447286 357368
rect 449898 357312 449954 357368
rect 451462 357312 451518 357368
rect 452658 357312 452714 357368
rect 454682 357312 454738 357368
rect 457534 357312 457590 357368
rect 462318 357312 462374 357368
rect 464342 357312 464398 357368
rect 467838 357312 467894 357368
rect 472622 357312 472678 357368
rect 477498 357312 477554 357368
rect 485778 357312 485834 357368
rect 433430 357176 433486 357232
rect 434626 357196 434682 357232
rect 434626 357176 434628 357196
rect 434628 357176 434680 357196
rect 434680 357176 434682 357196
rect 436006 357176 436062 357232
rect 438398 357176 438454 357232
rect 443090 357176 443146 357232
rect 441710 356516 441766 356552
rect 441710 356496 441712 356516
rect 441712 356496 441764 356516
rect 441764 356496 441766 356516
rect 442998 356496 443054 356552
rect 441986 356360 442042 356416
rect 445666 357076 445668 357096
rect 445668 357076 445720 357096
rect 445720 357076 445722 357096
rect 445666 357040 445722 357076
rect 445758 356632 445814 356688
rect 444378 356360 444434 356416
rect 447138 357040 447194 357096
rect 448518 356768 448574 356824
rect 448518 356496 448574 356552
rect 449990 357060 450046 357096
rect 449990 357040 449992 357060
rect 449992 357040 450044 357060
rect 450044 357040 450046 357060
rect 454038 357040 454094 357096
rect 452750 356924 452806 356960
rect 452750 356904 452752 356924
rect 452752 356904 452804 356924
rect 452804 356904 452806 356924
rect 456798 357212 456800 357232
rect 456800 357212 456852 357232
rect 456852 357212 456854 357232
rect 456798 357176 456854 357212
rect 455418 356904 455474 356960
rect 456798 356788 456854 356824
rect 456798 356768 456800 356788
rect 456800 356768 456852 356788
rect 456852 356768 456854 356788
rect 458178 357176 458234 357232
rect 460938 356108 460994 356144
rect 460938 356088 460940 356108
rect 460940 356088 460992 356108
rect 460992 356088 460994 356108
rect 470782 356224 470838 356280
rect 480534 357040 480590 357096
rect 474738 356360 474794 356416
rect 483018 356496 483074 356552
rect 498198 357312 498254 357368
rect 489918 356244 489974 356280
rect 489918 356224 489920 356244
rect 489920 356224 489972 356244
rect 489972 356224 489974 356244
rect 502338 356768 502394 356824
rect 500958 356360 501014 356416
rect 492678 356108 492734 356144
rect 492678 356088 492680 356108
rect 492680 356088 492732 356108
rect 492732 356088 492734 356108
rect 495438 356224 495494 356280
rect 505098 356108 505154 356144
rect 505098 356088 505100 356108
rect 505100 356088 505152 356108
rect 505152 356088 505154 356108
rect 456062 281968 456118 282024
rect 469862 281832 469918 281888
rect 517518 287136 517574 287192
rect 491942 281696 491998 281752
rect 514758 281560 514814 281616
rect 498934 233824 498990 233880
rect 538218 559136 538274 559192
rect 538218 439728 538274 439784
rect 542358 290536 542414 290592
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 617480 580226 617536
rect 579618 590960 579674 591016
rect 579618 577632 579674 577688
rect 579894 564304 579950 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579802 365064 579858 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580354 630808 580410 630864
rect 580446 418240 580502 418296
rect 580354 353912 580410 353968
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 548522 290400 548578 290456
rect 544382 284824 544438 284880
rect 513286 232464 513342 232520
rect 534814 230560 534870 230616
rect 532422 229200 532478 229256
rect 540334 280200 540390 280256
rect 580262 280880 580318 280936
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 205672 580226 205728
rect 580170 165824 580226 165880
rect 579802 139340 579804 139360
rect 579804 139340 579856 139360
rect 579856 139340 579858 139360
rect 579802 139304 579858 139340
rect 580170 125976 580226 126032
rect 579618 112784 579674 112840
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580446 280744 580502 280800
rect 580354 152632 580410 152688
rect 580722 219000 580778 219056
rect 580630 192480 580686 192536
rect 580538 179152 580594 179208
rect 580446 99456 580502 99512
rect 580262 59608 580318 59664
rect 580170 46280 580226 46336
rect 579986 19760 580042 19816
rect 579986 7520 580042 7576
rect 579986 6568 580042 6624
<< metal3 >>
rect 214414 700708 214420 700772
rect 214484 700770 214490 700772
rect 235165 700770 235231 700773
rect 214484 700768 235231 700770
rect 214484 700712 235170 700768
rect 235226 700712 235231 700768
rect 214484 700710 235231 700712
rect 214484 700708 214490 700710
rect 235165 700707 235231 700710
rect 211654 700572 211660 700636
rect 211724 700634 211730 700636
rect 267641 700634 267707 700637
rect 211724 700632 267707 700634
rect 211724 700576 267646 700632
rect 267702 700576 267707 700632
rect 211724 700574 267707 700576
rect 211724 700572 211730 700574
rect 267641 700571 267707 700574
rect 215886 700436 215892 700500
rect 215956 700498 215962 700500
rect 300117 700498 300183 700501
rect 215956 700496 300183 700498
rect 215956 700440 300122 700496
rect 300178 700440 300183 700496
rect 215956 700438 300183 700440
rect 215956 700436 215962 700438
rect 300117 700435 300183 700438
rect 395286 700436 395292 700500
rect 395356 700498 395362 700500
rect 494789 700498 494855 700501
rect 395356 700496 494855 700498
rect 395356 700440 494794 700496
rect 494850 700440 494855 700496
rect 395356 700438 494855 700440
rect 395356 700436 395362 700438
rect 494789 700435 494855 700438
rect 213126 700300 213132 700364
rect 213196 700362 213202 700364
rect 332501 700362 332567 700365
rect 213196 700360 332567 700362
rect 213196 700304 332506 700360
rect 332562 700304 332567 700360
rect 213196 700302 332567 700304
rect 213196 700300 213202 700302
rect 332501 700299 332567 700302
rect 398598 700300 398604 700364
rect 398668 700362 398674 700364
rect 527173 700362 527239 700365
rect 398668 700360 527239 700362
rect 398668 700304 527178 700360
rect 527234 700304 527239 700360
rect 398668 700302 527239 700304
rect 398668 700300 398674 700302
rect 527173 700299 527239 700302
rect 397453 699820 397519 699821
rect 397453 699818 397500 699820
rect 397408 699816 397500 699818
rect 397408 699760 397458 699816
rect 397408 699758 397500 699760
rect 397453 699756 397500 699758
rect 397564 699756 397570 699820
rect 397453 699755 397519 699756
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 170857 685948 170923 685949
rect 350993 685948 351059 685949
rect 530945 685948 531011 685949
rect 170806 685946 170812 685948
rect 170766 685886 170812 685946
rect 170876 685944 170923 685948
rect 350942 685946 350948 685948
rect 170918 685888 170923 685944
rect 170806 685884 170812 685886
rect 170876 685884 170923 685888
rect 350902 685886 350948 685946
rect 351012 685944 351059 685948
rect 530894 685946 530900 685948
rect 351054 685888 351059 685944
rect 350942 685884 350948 685886
rect 351012 685884 351059 685888
rect 530854 685886 530900 685946
rect 530964 685944 531011 685948
rect 531006 685888 531011 685944
rect 530894 685884 530900 685886
rect 530964 685884 531011 685888
rect 170857 685883 170923 685884
rect 350993 685883 351059 685884
rect 530945 685883 531011 685884
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect 176548 679160 177130 679220
rect 177070 679146 177130 679160
rect 178493 679146 178559 679149
rect 177070 679144 178559 679146
rect 177070 679088 178498 679144
rect 178554 679088 178559 679144
rect 177070 679086 178559 679088
rect 178493 679083 178559 679086
rect 356562 679010 356622 679190
rect 358813 679010 358879 679013
rect 356562 679008 358879 679010
rect 356562 678952 358818 679008
rect 358874 678952 358879 679008
rect 356562 678950 358879 678952
rect 536558 679010 536618 679190
rect 538213 679010 538279 679013
rect 536558 679008 538279 679010
rect 536558 678952 538218 679008
rect 538274 678952 538279 679008
rect 536558 678950 538279 678952
rect 358813 678947 358879 678950
rect 538213 678947 538279 678950
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 37825 636306 37891 636309
rect 39990 636306 40050 636894
rect 219390 636864 220064 636924
rect 399342 636864 400016 636924
rect 217225 636850 217291 636853
rect 219390 636850 219450 636864
rect 217225 636848 219450 636850
rect 217225 636792 217230 636848
rect 217286 636792 219450 636848
rect 217225 636790 219450 636792
rect 397269 636850 397335 636853
rect 399342 636850 399402 636864
rect 397269 636848 399402 636850
rect 397269 636792 397274 636848
rect 397330 636792 399402 636848
rect 397269 636790 399402 636792
rect 217225 636787 217291 636790
rect 397269 636787 397335 636790
rect 37825 636304 40050 636306
rect 37825 636248 37830 636304
rect 37886 636248 40050 636304
rect 37825 636246 40050 636248
rect 37825 636243 37891 636246
rect 38469 635354 38535 635357
rect 39990 635354 40050 635942
rect 219390 635912 220064 635972
rect 399342 635912 400016 635972
rect 217133 635898 217199 635901
rect 219390 635898 219450 635912
rect 217133 635896 219450 635898
rect 217133 635840 217138 635896
rect 217194 635840 219450 635896
rect 217133 635838 219450 635840
rect 396901 635898 396967 635901
rect 399342 635898 399402 635912
rect 396901 635896 399402 635898
rect 396901 635840 396906 635896
rect 396962 635840 399402 635896
rect 396901 635838 399402 635840
rect 217133 635835 217199 635838
rect 396901 635835 396967 635838
rect 38469 635352 40050 635354
rect 38469 635296 38474 635352
rect 38530 635296 40050 635352
rect 38469 635294 40050 635296
rect 38469 635291 38535 635294
rect 38510 633388 38516 633452
rect 38580 633450 38586 633452
rect 39990 633450 40050 633766
rect 219390 633736 220064 633796
rect 399342 633736 400016 633796
rect 217869 633722 217935 633725
rect 219390 633722 219450 633736
rect 217869 633720 219450 633722
rect 217869 633664 217874 633720
rect 217930 633664 219450 633720
rect 217869 633662 219450 633664
rect 396993 633722 397059 633725
rect 399342 633722 399402 633736
rect 396993 633720 399402 633722
rect 396993 633664 396998 633720
rect 397054 633664 399402 633720
rect 396993 633662 399402 633664
rect 217869 633659 217935 633662
rect 396993 633659 397059 633662
rect 38580 633390 40050 633450
rect 38580 633388 38586 633390
rect 38009 632226 38075 632229
rect 39990 632226 40050 632814
rect 219390 632784 220064 632844
rect 399342 632784 400016 632844
rect 217685 632770 217751 632773
rect 219390 632770 219450 632784
rect 217685 632768 219450 632770
rect 217685 632712 217690 632768
rect 217746 632712 219450 632768
rect 217685 632710 219450 632712
rect 396625 632770 396691 632773
rect 399342 632770 399402 632784
rect 396625 632768 399402 632770
rect 396625 632712 396630 632768
rect 396686 632712 399402 632768
rect 396625 632710 399402 632712
rect 217685 632707 217751 632710
rect 396625 632707 396691 632710
rect 38009 632224 40050 632226
rect -960 632090 480 632180
rect 38009 632168 38014 632224
rect 38070 632168 40050 632224
rect 38009 632166 40050 632168
rect 38009 632163 38075 632166
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 38101 630730 38167 630733
rect 39990 630730 40050 631046
rect 219390 631016 220064 631076
rect 399342 631016 400016 631076
rect 217593 631002 217659 631005
rect 219390 631002 219450 631016
rect 217593 631000 219450 631002
rect 217593 630944 217598 631000
rect 217654 630944 219450 631000
rect 217593 630942 219450 630944
rect 397085 631002 397151 631005
rect 399342 631002 399402 631016
rect 397085 631000 399402 631002
rect 397085 630944 397090 631000
rect 397146 630944 399402 631000
rect 397085 630942 399402 630944
rect 217593 630939 217659 630942
rect 397085 630939 397151 630942
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 38101 630728 40050 630730
rect 38101 630672 38106 630728
rect 38162 630672 40050 630728
rect 583520 630716 584960 630806
rect 38101 630670 40050 630672
rect 38101 630667 38167 630670
rect 38285 629370 38351 629373
rect 39990 629370 40050 629958
rect 219390 629928 220064 629988
rect 399342 629928 400016 629988
rect 217501 629914 217567 629917
rect 219390 629914 219450 629928
rect 217501 629912 219450 629914
rect 217501 629856 217506 629912
rect 217562 629856 219450 629912
rect 217501 629854 219450 629856
rect 397361 629914 397427 629917
rect 399342 629914 399402 629928
rect 397361 629912 399402 629914
rect 397361 629856 397366 629912
rect 397422 629856 399402 629912
rect 397361 629854 399402 629856
rect 217501 629851 217567 629854
rect 397361 629851 397427 629854
rect 38285 629368 40050 629370
rect 38285 629312 38290 629368
rect 38346 629312 40050 629368
rect 38285 629310 40050 629312
rect 38285 629307 38351 629310
rect 38193 628010 38259 628013
rect 39990 628010 40050 628190
rect 219390 628160 220064 628220
rect 399342 628160 400016 628220
rect 217409 628146 217475 628149
rect 219390 628146 219450 628160
rect 217409 628144 219450 628146
rect 217409 628088 217414 628144
rect 217470 628088 219450 628144
rect 217409 628086 219450 628088
rect 396809 628146 396875 628149
rect 399342 628146 399402 628160
rect 396809 628144 399402 628146
rect 396809 628088 396814 628144
rect 396870 628088 399402 628144
rect 396809 628086 399402 628088
rect 217409 628083 217475 628086
rect 396809 628083 396875 628086
rect 38193 628008 40050 628010
rect 38193 627952 38198 628008
rect 38254 627952 40050 628008
rect 38193 627950 40050 627952
rect 38193 627947 38259 627950
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 38561 610058 38627 610061
rect 217777 610058 217843 610061
rect 396717 610058 396783 610061
rect 38561 610056 40050 610058
rect 38561 610000 38566 610056
rect 38622 610000 40050 610056
rect 38561 609998 40050 610000
rect 38561 609995 38627 609998
rect 39990 609966 40050 609998
rect 217777 610056 219450 610058
rect 217777 610000 217782 610056
rect 217838 610000 219450 610056
rect 217777 609998 219450 610000
rect 217777 609995 217843 609998
rect 219390 609996 219450 609998
rect 396717 610056 399402 610058
rect 396717 610000 396722 610056
rect 396778 610000 399402 610056
rect 396717 609998 399402 610000
rect 219390 609936 220064 609996
rect 396717 609995 396783 609998
rect 399342 609996 399402 609998
rect 399342 609936 400016 609996
rect 38326 608364 38332 608428
rect 38396 608426 38402 608428
rect 38396 608366 40050 608426
rect 38396 608364 38402 608366
rect 39990 608334 40050 608366
rect 219390 608304 220064 608364
rect 399342 608304 400016 608364
rect 216673 608290 216739 608293
rect 219390 608290 219450 608304
rect 216673 608288 219450 608290
rect 216673 608232 216678 608288
rect 216734 608232 219450 608288
rect 216673 608230 219450 608232
rect 397177 608290 397243 608293
rect 399342 608290 399402 608304
rect 397177 608288 399402 608290
rect 397177 608232 397182 608288
rect 397238 608232 399402 608288
rect 397177 608230 399402 608232
rect 216673 608227 216739 608230
rect 397177 608227 397243 608230
rect 38694 607412 38700 607476
rect 38764 607474 38770 607476
rect 39990 607474 40050 608062
rect 219390 608032 220064 608092
rect 399342 608032 400016 608092
rect 219198 607956 219204 608020
rect 219268 608018 219274 608020
rect 219390 608018 219450 608032
rect 219268 607958 219450 608018
rect 219268 607956 219274 607958
rect 38764 607414 40050 607474
rect 38764 607412 38770 607414
rect 357934 607412 357940 607476
rect 358004 607474 358010 607476
rect 399342 607474 399402 608032
rect 358004 607414 399402 607474
rect 358004 607412 358010 607414
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect 258073 599588 258139 599589
rect 258073 599584 258086 599588
rect 258150 599586 258156 599588
rect 277301 599586 277367 599589
rect 435909 599588 435975 599589
rect 278480 599586 278486 599588
rect 258073 599528 258078 599584
rect 258073 599524 258086 599528
rect 258150 599526 258230 599586
rect 277301 599584 278486 599586
rect 277301 599528 277306 599584
rect 277362 599528 278486 599584
rect 277301 599526 278486 599528
rect 258150 599524 258156 599526
rect 258073 599523 258139 599524
rect 277301 599523 277367 599526
rect 278480 599524 278486 599526
rect 278550 599524 278556 599588
rect 435904 599586 435910 599588
rect 435818 599526 435910 599586
rect 435904 599524 435910 599526
rect 435974 599524 435980 599588
rect 450854 599524 450860 599588
rect 450924 599586 450930 599588
rect 451136 599586 451142 599588
rect 450924 599526 451142 599586
rect 450924 599524 450930 599526
rect 451136 599524 451142 599526
rect 451206 599524 451212 599588
rect 435909 599523 435975 599524
rect 451089 599450 451155 599453
rect 452142 599450 452148 599452
rect 451089 599448 452148 599450
rect 451089 599392 451094 599448
rect 451150 599392 452148 599448
rect 451089 599390 452148 599392
rect 451089 599387 451155 599390
rect 452142 599388 452148 599390
rect 452212 599388 452218 599452
rect 56409 597546 56475 597549
rect 63217 597548 63283 597549
rect 61694 597546 61700 597548
rect 56409 597544 61700 597546
rect 56409 597488 56414 597544
rect 56470 597488 61700 597544
rect 56409 597486 61700 597488
rect 56409 597483 56475 597486
rect 61694 597484 61700 597486
rect 61764 597484 61770 597548
rect 63166 597546 63172 597548
rect 63126 597486 63172 597546
rect 63236 597544 63283 597548
rect 63278 597488 63283 597544
rect 63166 597484 63172 597486
rect 63236 597484 63283 597488
rect 63217 597483 63283 597484
rect 64229 597548 64295 597549
rect 64229 597544 64276 597548
rect 64340 597546 64346 597548
rect 64229 597488 64234 597544
rect 64229 597484 64276 597488
rect 64340 597486 64386 597546
rect 64340 597484 64346 597486
rect 64638 597484 64644 597548
rect 64708 597546 64714 597548
rect 64873 597546 64939 597549
rect 64708 597544 64939 597546
rect 64708 597488 64878 597544
rect 64934 597488 64939 597544
rect 64708 597486 64939 597488
rect 64708 597484 64714 597486
rect 64229 597483 64295 597484
rect 64873 597483 64939 597486
rect 66478 597484 66484 597548
rect 66548 597546 66554 597548
rect 66805 597546 66871 597549
rect 67633 597548 67699 597549
rect 67582 597546 67588 597548
rect 66548 597544 66871 597546
rect 66548 597488 66810 597544
rect 66866 597488 66871 597544
rect 66548 597486 66871 597488
rect 67542 597486 67588 597546
rect 67652 597544 67699 597548
rect 67694 597488 67699 597544
rect 66548 597484 66554 597486
rect 66805 597483 66871 597486
rect 67582 597484 67588 597486
rect 67652 597484 67699 597488
rect 68318 597484 68324 597548
rect 68388 597546 68394 597548
rect 68921 597546 68987 597549
rect 68388 597544 68987 597546
rect 68388 597488 68926 597544
rect 68982 597488 68987 597544
rect 68388 597486 68987 597488
rect 68388 597484 68394 597486
rect 67633 597483 67699 597484
rect 68921 597483 68987 597486
rect 69749 597546 69815 597549
rect 69974 597546 69980 597548
rect 69749 597544 69980 597546
rect 69749 597488 69754 597544
rect 69810 597488 69980 597544
rect 69749 597486 69980 597488
rect 69749 597483 69815 597486
rect 69974 597484 69980 597486
rect 70044 597484 70050 597548
rect 70710 597484 70716 597548
rect 70780 597546 70786 597548
rect 71681 597546 71747 597549
rect 70780 597544 71747 597546
rect 70780 597488 71686 597544
rect 71742 597488 71747 597544
rect 70780 597486 71747 597488
rect 70780 597484 70786 597486
rect 71681 597483 71747 597486
rect 73153 597546 73219 597549
rect 73470 597546 73476 597548
rect 73153 597544 73476 597546
rect 73153 597488 73158 597544
rect 73214 597488 73476 597544
rect 73153 597486 73476 597488
rect 73153 597483 73219 597486
rect 73470 597484 73476 597486
rect 73540 597484 73546 597548
rect 73654 597484 73660 597548
rect 73724 597546 73730 597548
rect 74441 597546 74507 597549
rect 73724 597544 74507 597546
rect 73724 597488 74446 597544
rect 74502 597488 74507 597544
rect 73724 597486 74507 597488
rect 73724 597484 73730 597486
rect 74441 597483 74507 597486
rect 74574 597484 74580 597548
rect 74644 597546 74650 597548
rect 74901 597546 74967 597549
rect 74644 597544 74967 597546
rect 74644 597488 74906 597544
rect 74962 597488 74967 597544
rect 74644 597486 74967 597488
rect 74644 597484 74650 597486
rect 74901 597483 74967 597486
rect 76046 597484 76052 597548
rect 76116 597546 76122 597548
rect 77201 597546 77267 597549
rect 76116 597544 77267 597546
rect 76116 597488 77206 597544
rect 77262 597488 77267 597544
rect 76116 597486 77267 597488
rect 76116 597484 76122 597486
rect 77201 597483 77267 597486
rect 78029 597548 78095 597549
rect 78029 597544 78076 597548
rect 78140 597546 78146 597548
rect 78029 597488 78034 597544
rect 78029 597484 78076 597488
rect 78140 597486 78186 597546
rect 78140 597484 78146 597486
rect 78438 597484 78444 597548
rect 78508 597546 78514 597548
rect 78581 597546 78647 597549
rect 78508 597544 78647 597546
rect 78508 597488 78586 597544
rect 78642 597488 78647 597544
rect 78508 597486 78647 597488
rect 78508 597484 78514 597486
rect 78029 597483 78095 597484
rect 78581 597483 78647 597486
rect 81014 597484 81020 597548
rect 81084 597546 81090 597548
rect 81341 597546 81407 597549
rect 81084 597544 81407 597546
rect 81084 597488 81346 597544
rect 81402 597488 81407 597544
rect 81084 597486 81407 597488
rect 81084 597484 81090 597486
rect 81341 597483 81407 597486
rect 83958 597484 83964 597548
rect 84028 597546 84034 597548
rect 84193 597546 84259 597549
rect 84028 597544 84259 597546
rect 84028 597488 84198 597544
rect 84254 597488 84259 597544
rect 84028 597486 84259 597488
rect 84028 597484 84034 597486
rect 84193 597483 84259 597486
rect 85982 597484 85988 597548
rect 86052 597546 86058 597548
rect 86861 597546 86927 597549
rect 88241 597548 88307 597549
rect 86052 597544 86927 597546
rect 86052 597488 86866 597544
rect 86922 597488 86927 597544
rect 86052 597486 86927 597488
rect 86052 597484 86058 597486
rect 86861 597483 86927 597486
rect 88190 597484 88196 597548
rect 88260 597546 88307 597548
rect 92473 597546 92539 597549
rect 93342 597546 93348 597548
rect 88260 597544 88352 597546
rect 88302 597488 88352 597544
rect 88260 597486 88352 597488
rect 92473 597544 93348 597546
rect 92473 597488 92478 597544
rect 92534 597488 93348 597544
rect 92473 597486 93348 597488
rect 88260 597484 88307 597486
rect 88241 597483 88307 597484
rect 92473 597483 92539 597486
rect 93342 597484 93348 597486
rect 93412 597484 93418 597548
rect 93526 597484 93532 597548
rect 93596 597546 93602 597548
rect 93761 597546 93827 597549
rect 93596 597544 93827 597546
rect 93596 597488 93766 597544
rect 93822 597488 93827 597544
rect 93596 597486 93827 597488
rect 93596 597484 93602 597486
rect 93761 597483 93827 597486
rect 122598 597484 122604 597548
rect 122668 597546 122674 597548
rect 124121 597546 124187 597549
rect 122668 597544 124187 597546
rect 122668 597488 124126 597544
rect 124182 597488 124187 597544
rect 122668 597486 124187 597488
rect 122668 597484 122674 597486
rect 124121 597483 124187 597486
rect 128486 597484 128492 597548
rect 128556 597546 128562 597548
rect 129641 597546 129707 597549
rect 131021 597548 131087 597549
rect 131021 597546 131068 597548
rect 128556 597544 129707 597546
rect 128556 597488 129646 597544
rect 129702 597488 129707 597544
rect 128556 597486 129707 597488
rect 130976 597544 131068 597546
rect 130976 597488 131026 597544
rect 130976 597486 131068 597488
rect 128556 597484 128562 597486
rect 129641 597483 129707 597486
rect 131021 597484 131068 597486
rect 131132 597484 131138 597548
rect 133454 597484 133460 597548
rect 133524 597546 133530 597548
rect 133781 597546 133847 597549
rect 133524 597544 133847 597546
rect 133524 597488 133786 597544
rect 133842 597488 133847 597544
rect 133524 597486 133847 597488
rect 133524 597484 133530 597486
rect 131021 597483 131087 597484
rect 133781 597483 133847 597486
rect 135846 597484 135852 597548
rect 135916 597546 135922 597548
rect 136541 597546 136607 597549
rect 135916 597544 136607 597546
rect 135916 597488 136546 597544
rect 136602 597488 136607 597544
rect 135916 597486 136607 597488
rect 135916 597484 135922 597486
rect 136541 597483 136607 597486
rect 140998 597484 141004 597548
rect 141068 597546 141074 597548
rect 142061 597546 142127 597549
rect 141068 597544 142127 597546
rect 141068 597488 142066 597544
rect 142122 597488 142127 597544
rect 141068 597486 142127 597488
rect 141068 597484 141074 597486
rect 142061 597483 142127 597486
rect 145966 597484 145972 597548
rect 146036 597546 146042 597548
rect 146201 597546 146267 597549
rect 235993 597548 236059 597549
rect 146036 597544 146267 597546
rect 146036 597488 146206 597544
rect 146262 597488 146267 597544
rect 146036 597486 146267 597488
rect 146036 597484 146042 597486
rect 146201 597483 146267 597486
rect 235942 597484 235948 597548
rect 236012 597546 236059 597548
rect 236177 597546 236243 597549
rect 237046 597546 237052 597548
rect 236012 597544 236104 597546
rect 236054 597488 236104 597544
rect 236012 597486 236104 597488
rect 236177 597544 237052 597546
rect 236177 597488 236182 597544
rect 236238 597488 237052 597544
rect 236177 597486 237052 597488
rect 236012 597484 236059 597486
rect 235993 597483 236059 597484
rect 236177 597483 236243 597486
rect 237046 597484 237052 597486
rect 237116 597484 237122 597548
rect 237373 597546 237439 597549
rect 243077 597548 243143 597549
rect 244273 597548 244339 597549
rect 238150 597546 238156 597548
rect 237373 597544 238156 597546
rect 237373 597488 237378 597544
rect 237434 597488 238156 597544
rect 237373 597486 238156 597488
rect 237373 597483 237439 597486
rect 238150 597484 238156 597486
rect 238220 597484 238226 597548
rect 243077 597544 243124 597548
rect 243188 597546 243194 597548
rect 244222 597546 244228 597548
rect 243077 597488 243082 597544
rect 243077 597484 243124 597488
rect 243188 597486 243234 597546
rect 244182 597486 244228 597546
rect 244292 597544 244339 597548
rect 244334 597488 244339 597544
rect 243188 597484 243194 597486
rect 244222 597484 244228 597486
rect 244292 597484 244339 597488
rect 243077 597483 243143 597484
rect 244273 597483 244339 597484
rect 245469 597548 245535 597549
rect 246481 597548 246547 597549
rect 245469 597544 245516 597548
rect 245580 597546 245586 597548
rect 246430 597546 246436 597548
rect 245469 597488 245474 597544
rect 245469 597484 245516 597488
rect 245580 597486 245626 597546
rect 246390 597486 246436 597546
rect 246500 597544 246547 597548
rect 246542 597488 246547 597544
rect 245580 597484 245586 597486
rect 246430 597484 246436 597486
rect 246500 597484 246547 597488
rect 245469 597483 245535 597484
rect 246481 597483 246547 597484
rect 247033 597546 247099 597549
rect 248270 597546 248276 597548
rect 247033 597544 248276 597546
rect 247033 597488 247038 597544
rect 247094 597488 248276 597544
rect 247033 597486 248276 597488
rect 247033 597483 247099 597486
rect 248270 597484 248276 597486
rect 248340 597484 248346 597548
rect 248413 597546 248479 597549
rect 248638 597546 248644 597548
rect 248413 597544 248644 597546
rect 248413 597488 248418 597544
rect 248474 597488 248644 597544
rect 248413 597486 248644 597488
rect 248413 597483 248479 597486
rect 248638 597484 248644 597486
rect 248708 597484 248714 597548
rect 249793 597546 249859 597549
rect 250662 597546 250668 597548
rect 249793 597544 250668 597546
rect 249793 597488 249798 597544
rect 249854 597488 250668 597544
rect 249793 597486 250668 597488
rect 249793 597483 249859 597486
rect 250662 597484 250668 597486
rect 250732 597484 250738 597548
rect 252093 597546 252159 597549
rect 253473 597548 253539 597549
rect 254577 597548 254643 597549
rect 252318 597546 252324 597548
rect 252093 597544 252324 597546
rect 252093 597488 252098 597544
rect 252154 597488 252324 597544
rect 252093 597486 252324 597488
rect 252093 597483 252159 597486
rect 252318 597484 252324 597486
rect 252388 597484 252394 597548
rect 253422 597484 253428 597548
rect 253492 597546 253539 597548
rect 254526 597546 254532 597548
rect 253492 597544 253584 597546
rect 253534 597488 253584 597544
rect 253492 597486 253584 597488
rect 254486 597486 254532 597546
rect 254596 597544 254643 597548
rect 254638 597488 254643 597544
rect 253492 597484 253539 597486
rect 254526 597484 254532 597486
rect 254596 597484 254643 597488
rect 253473 597483 253539 597484
rect 254577 597483 254643 597484
rect 255405 597546 255471 597549
rect 255814 597546 255820 597548
rect 255405 597544 255820 597546
rect 255405 597488 255410 597544
rect 255466 597488 255820 597544
rect 255405 597486 255820 597488
rect 255405 597483 255471 597486
rect 255814 597484 255820 597486
rect 255884 597484 255890 597548
rect 256693 597546 256759 597549
rect 256918 597546 256924 597548
rect 256693 597544 256924 597546
rect 256693 597488 256698 597544
rect 256754 597488 256924 597544
rect 256693 597486 256924 597488
rect 256693 597483 256759 597486
rect 256918 597484 256924 597486
rect 256988 597484 256994 597548
rect 260833 597546 260899 597549
rect 263593 597548 263659 597549
rect 261702 597546 261708 597548
rect 260833 597544 261708 597546
rect 260833 597488 260838 597544
rect 260894 597488 261708 597544
rect 260833 597486 261708 597488
rect 260833 597483 260899 597486
rect 261702 597484 261708 597486
rect 261772 597484 261778 597548
rect 263542 597484 263548 597548
rect 263612 597546 263659 597548
rect 264973 597546 265039 597549
rect 265934 597546 265940 597548
rect 263612 597544 263704 597546
rect 263654 597488 263704 597544
rect 263612 597486 263704 597488
rect 264973 597544 265940 597546
rect 264973 597488 264978 597544
rect 265034 597488 265940 597544
rect 264973 597486 265940 597488
rect 263612 597484 263659 597486
rect 263593 597483 263659 597484
rect 264973 597483 265039 597486
rect 265934 597484 265940 597486
rect 266004 597484 266010 597548
rect 267733 597546 267799 597549
rect 268326 597546 268332 597548
rect 267733 597544 268332 597546
rect 267733 597488 267738 597544
rect 267794 597488 268332 597544
rect 267733 597486 268332 597488
rect 267733 597483 267799 597486
rect 268326 597484 268332 597486
rect 268396 597484 268402 597548
rect 270493 597546 270559 597549
rect 270902 597546 270908 597548
rect 270493 597544 270908 597546
rect 270493 597488 270498 597544
rect 270554 597488 270908 597544
rect 270493 597486 270908 597488
rect 270493 597483 270559 597486
rect 270902 597484 270908 597486
rect 270972 597484 270978 597548
rect 276013 597546 276079 597549
rect 276974 597546 276980 597548
rect 276013 597544 276980 597546
rect 276013 597488 276018 597544
rect 276074 597488 276980 597544
rect 276013 597486 276980 597488
rect 276013 597483 276079 597486
rect 276974 597484 276980 597486
rect 277044 597484 277050 597548
rect 280153 597546 280219 597549
rect 280838 597546 280844 597548
rect 280153 597544 280844 597546
rect 280153 597488 280158 597544
rect 280214 597488 280844 597544
rect 280153 597486 280844 597488
rect 280153 597483 280219 597486
rect 280838 597484 280844 597486
rect 280908 597484 280914 597548
rect 282913 597546 282979 597549
rect 283414 597546 283420 597548
rect 282913 597544 283420 597546
rect 282913 597488 282918 597544
rect 282974 597488 283420 597544
rect 282913 597486 283420 597488
rect 282913 597483 282979 597486
rect 283414 597484 283420 597486
rect 283484 597484 283490 597548
rect 285673 597546 285739 597549
rect 285990 597546 285996 597548
rect 285673 597544 285996 597546
rect 285673 597488 285678 597544
rect 285734 597488 285996 597544
rect 285673 597486 285996 597488
rect 285673 597483 285739 597486
rect 285990 597484 285996 597486
rect 286060 597484 286066 597548
rect 289813 597546 289879 597549
rect 290958 597546 290964 597548
rect 289813 597544 290964 597546
rect 289813 597488 289818 597544
rect 289874 597488 290964 597544
rect 289813 597486 290964 597488
rect 289813 597483 289879 597486
rect 290958 597484 290964 597486
rect 291028 597484 291034 597548
rect 292573 597546 292639 597549
rect 293350 597546 293356 597548
rect 292573 597544 293356 597546
rect 292573 597488 292578 597544
rect 292634 597488 293356 597544
rect 292573 597486 293356 597488
rect 292573 597483 292639 597486
rect 293350 597484 293356 597486
rect 293420 597484 293426 597548
rect 415393 597546 415459 597549
rect 416078 597546 416084 597548
rect 415393 597544 416084 597546
rect 415393 597488 415398 597544
rect 415454 597488 416084 597544
rect 415393 597486 416084 597488
rect 415393 597483 415459 597486
rect 416078 597484 416084 597486
rect 416148 597484 416154 597548
rect 416773 597546 416839 597549
rect 417182 597546 417188 597548
rect 416773 597544 417188 597546
rect 416773 597488 416778 597544
rect 416834 597488 417188 597544
rect 416773 597486 417188 597488
rect 416773 597483 416839 597486
rect 417182 597484 417188 597486
rect 417252 597484 417258 597548
rect 418153 597546 418219 597549
rect 418286 597546 418292 597548
rect 418153 597544 418292 597546
rect 418153 597488 418158 597544
rect 418214 597488 418292 597544
rect 418153 597486 418292 597488
rect 418153 597483 418219 597486
rect 418286 597484 418292 597486
rect 418356 597484 418362 597548
rect 419533 597546 419599 597549
rect 420494 597546 420500 597548
rect 419533 597544 420500 597546
rect 419533 597488 419538 597544
rect 419594 597488 420500 597544
rect 419533 597486 420500 597488
rect 419533 597483 419599 597486
rect 420494 597484 420500 597486
rect 420564 597484 420570 597548
rect 420913 597546 420979 597549
rect 423121 597548 423187 597549
rect 421782 597546 421788 597548
rect 420913 597544 421788 597546
rect 420913 597488 420918 597544
rect 420974 597488 421788 597544
rect 420913 597486 421788 597488
rect 420913 597483 420979 597486
rect 421782 597484 421788 597486
rect 421852 597484 421858 597548
rect 423070 597546 423076 597548
rect 423030 597486 423076 597546
rect 423140 597544 423187 597548
rect 423182 597488 423187 597544
rect 423070 597484 423076 597486
rect 423140 597484 423187 597488
rect 424174 597484 424180 597548
rect 424244 597546 424250 597548
rect 424961 597546 425027 597549
rect 424244 597544 425027 597546
rect 424244 597488 424966 597544
rect 425022 597488 425027 597544
rect 424244 597486 425027 597488
rect 424244 597484 424250 597486
rect 423121 597483 423187 597484
rect 424961 597483 425027 597486
rect 425462 597484 425468 597548
rect 425532 597546 425538 597548
rect 425605 597546 425671 597549
rect 425532 597544 425671 597546
rect 425532 597488 425610 597544
rect 425666 597488 425671 597544
rect 425532 597486 425671 597488
rect 425532 597484 425538 597486
rect 425605 597483 425671 597486
rect 426525 597548 426591 597549
rect 427629 597548 427695 597549
rect 426525 597544 426572 597548
rect 426636 597546 426642 597548
rect 426525 597488 426530 597544
rect 426525 597484 426572 597488
rect 426636 597486 426682 597546
rect 427629 597544 427676 597548
rect 427740 597546 427746 597548
rect 427997 597546 428063 597549
rect 428590 597546 428596 597548
rect 427629 597488 427634 597544
rect 426636 597484 426642 597486
rect 427629 597484 427676 597488
rect 427740 597486 427786 597546
rect 427997 597544 428596 597546
rect 427997 597488 428002 597544
rect 428058 597488 428596 597544
rect 427997 597486 428596 597488
rect 427740 597484 427746 597486
rect 426525 597483 426591 597484
rect 427629 597483 427695 597484
rect 427997 597483 428063 597486
rect 428590 597484 428596 597486
rect 428660 597484 428666 597548
rect 429193 597546 429259 597549
rect 430573 597548 430639 597549
rect 430062 597546 430068 597548
rect 429193 597544 430068 597546
rect 429193 597488 429198 597544
rect 429254 597488 430068 597544
rect 429193 597486 430068 597488
rect 429193 597483 429259 597486
rect 430062 597484 430068 597486
rect 430132 597484 430138 597548
rect 430573 597546 430620 597548
rect 430528 597544 430620 597546
rect 430528 597488 430578 597544
rect 430528 597486 430620 597488
rect 430573 597484 430620 597486
rect 430684 597484 430690 597548
rect 433333 597546 433399 597549
rect 434529 597548 434595 597549
rect 433742 597546 433748 597548
rect 433333 597544 433748 597546
rect 433333 597488 433338 597544
rect 433394 597488 433748 597544
rect 433333 597486 433748 597488
rect 430573 597483 430639 597484
rect 433333 597483 433399 597486
rect 433742 597484 433748 597486
rect 433812 597484 433818 597548
rect 434478 597546 434484 597548
rect 434438 597486 434484 597546
rect 434548 597544 434595 597548
rect 434590 597488 434595 597544
rect 434478 597484 434484 597486
rect 434548 597484 434595 597488
rect 434529 597483 434595 597484
rect 434713 597546 434779 597549
rect 437105 597548 437171 597549
rect 435950 597546 435956 597548
rect 434713 597544 435956 597546
rect 434713 597488 434718 597544
rect 434774 597488 435956 597544
rect 434713 597486 435956 597488
rect 434713 597483 434779 597486
rect 435950 597484 435956 597486
rect 436020 597484 436026 597548
rect 437054 597546 437060 597548
rect 437014 597486 437060 597546
rect 437124 597544 437171 597548
rect 437166 597488 437171 597544
rect 437054 597484 437060 597486
rect 437124 597484 437171 597488
rect 437105 597483 437171 597484
rect 437473 597546 437539 597549
rect 437974 597546 437980 597548
rect 437473 597544 437980 597546
rect 437473 597488 437478 597544
rect 437534 597488 437980 597544
rect 437473 597486 437980 597488
rect 437473 597483 437539 597486
rect 437974 597484 437980 597486
rect 438044 597484 438050 597548
rect 438853 597546 438919 597549
rect 439446 597546 439452 597548
rect 438853 597544 439452 597546
rect 438853 597488 438858 597544
rect 438914 597488 439452 597544
rect 438853 597486 439452 597488
rect 438853 597483 438919 597486
rect 439446 597484 439452 597486
rect 439516 597484 439522 597548
rect 441981 597546 442047 597549
rect 442758 597546 442764 597548
rect 441981 597544 442764 597546
rect 441981 597488 441986 597544
rect 442042 597488 442764 597544
rect 441981 597486 442764 597488
rect 441981 597483 442047 597486
rect 442758 597484 442764 597486
rect 442828 597484 442834 597548
rect 442993 597546 443059 597549
rect 443494 597546 443500 597548
rect 442993 597544 443500 597546
rect 442993 597488 442998 597544
rect 443054 597488 443500 597544
rect 442993 597486 443500 597488
rect 442993 597483 443059 597486
rect 443494 597484 443500 597486
rect 443564 597484 443570 597548
rect 443637 597546 443703 597549
rect 443862 597546 443868 597548
rect 443637 597544 443868 597546
rect 443637 597488 443642 597544
rect 443698 597488 443868 597544
rect 443637 597486 443868 597488
rect 443637 597483 443703 597486
rect 443862 597484 443868 597486
rect 443932 597484 443938 597548
rect 444373 597546 444439 597549
rect 445334 597546 445340 597548
rect 444373 597544 445340 597546
rect 444373 597488 444378 597544
rect 444434 597488 445340 597544
rect 444373 597486 445340 597488
rect 444373 597483 444439 597486
rect 445334 597484 445340 597486
rect 445404 597484 445410 597548
rect 445753 597546 445819 597549
rect 445886 597546 445892 597548
rect 445753 597544 445892 597546
rect 445753 597488 445758 597544
rect 445814 597488 445892 597544
rect 445753 597486 445892 597488
rect 445753 597483 445819 597486
rect 445886 597484 445892 597486
rect 445956 597484 445962 597548
rect 447133 597546 447199 597549
rect 448278 597546 448284 597548
rect 447133 597544 448284 597546
rect 447133 597488 447138 597544
rect 447194 597488 448284 597544
rect 447133 597486 448284 597488
rect 447133 597483 447199 597486
rect 448278 597484 448284 597486
rect 448348 597484 448354 597548
rect 449893 597546 449959 597549
rect 451038 597546 451044 597548
rect 449893 597544 451044 597546
rect 449893 597488 449898 597544
rect 449954 597488 451044 597544
rect 449893 597486 451044 597488
rect 449893 597483 449959 597486
rect 451038 597484 451044 597486
rect 451108 597484 451114 597548
rect 456006 597546 456012 597548
rect 451230 597486 456012 597546
rect 39849 597410 39915 597413
rect 58198 597410 58204 597412
rect 39849 597408 58204 597410
rect 39849 597352 39854 597408
rect 39910 597352 58204 597408
rect 39849 597350 58204 597352
rect 39849 597347 39915 597350
rect 58198 597348 58204 597350
rect 58268 597348 58274 597412
rect 68686 597348 68692 597412
rect 68756 597410 68762 597412
rect 68829 597410 68895 597413
rect 71313 597412 71379 597413
rect 71262 597410 71268 597412
rect 68756 597408 68895 597410
rect 68756 597352 68834 597408
rect 68890 597352 68895 597408
rect 68756 597350 68895 597352
rect 71222 597350 71268 597410
rect 71332 597408 71379 597412
rect 71374 597352 71379 597408
rect 68756 597348 68762 597350
rect 68829 597347 68895 597350
rect 71262 597348 71268 597350
rect 71332 597348 71379 597352
rect 71313 597347 71379 597348
rect 71773 597410 71839 597413
rect 72366 597410 72372 597412
rect 71773 597408 72372 597410
rect 71773 597352 71778 597408
rect 71834 597352 72372 597408
rect 71773 597350 72372 597352
rect 71773 597347 71839 597350
rect 72366 597348 72372 597350
rect 72436 597348 72442 597412
rect 75862 597348 75868 597412
rect 75932 597410 75938 597412
rect 76005 597410 76071 597413
rect 75932 597408 76071 597410
rect 75932 597352 76010 597408
rect 76066 597352 76071 597408
rect 75932 597350 76071 597352
rect 75932 597348 75938 597350
rect 76005 597347 76071 597350
rect 76966 597348 76972 597412
rect 77036 597410 77042 597412
rect 77109 597410 77175 597413
rect 77036 597408 77175 597410
rect 77036 597352 77114 597408
rect 77170 597352 77175 597408
rect 77036 597350 77175 597352
rect 77036 597348 77042 597350
rect 77109 597347 77175 597350
rect 82813 597410 82879 597413
rect 83774 597410 83780 597412
rect 82813 597408 83780 597410
rect 82813 597352 82818 597408
rect 82874 597352 83780 597408
rect 82813 597350 83780 597352
rect 82813 597347 82879 597350
rect 83774 597348 83780 597350
rect 83844 597348 83850 597412
rect 98126 597410 98132 597412
rect 84150 597350 98132 597410
rect 39798 597212 39804 597276
rect 39868 597274 39874 597276
rect 60590 597274 60596 597276
rect 39868 597214 60596 597274
rect 39868 597212 39874 597214
rect 60590 597212 60596 597214
rect 60660 597212 60666 597276
rect 81433 597274 81499 597277
rect 81750 597274 81756 597276
rect 81433 597272 81756 597274
rect 81433 597216 81438 597272
rect 81494 597216 81756 597272
rect 81433 597214 81756 597216
rect 81433 597211 81499 597214
rect 81750 597212 81756 597214
rect 81820 597212 81826 597276
rect 39573 597138 39639 597141
rect 56409 597138 56475 597141
rect 39573 597136 56475 597138
rect 39573 597080 39578 597136
rect 39634 597080 56414 597136
rect 56470 597080 56475 597136
rect 39573 597078 56475 597080
rect 39573 597075 39639 597078
rect 56409 597075 56475 597078
rect 56593 597138 56659 597141
rect 57094 597138 57100 597140
rect 56593 597136 57100 597138
rect 56593 597080 56598 597136
rect 56654 597080 57100 597136
rect 56593 597078 57100 597080
rect 56593 597075 56659 597078
rect 57094 597076 57100 597078
rect 57164 597076 57170 597140
rect 59353 597138 59419 597141
rect 59486 597138 59492 597140
rect 59353 597136 59492 597138
rect 59353 597080 59358 597136
rect 59414 597080 59492 597136
rect 59353 597078 59492 597080
rect 59353 597075 59419 597078
rect 59486 597076 59492 597078
rect 59556 597076 59562 597140
rect 84150 597138 84210 597350
rect 98126 597348 98132 597350
rect 98196 597348 98202 597412
rect 108246 597348 108252 597412
rect 108316 597410 108322 597412
rect 108941 597410 109007 597413
rect 108316 597408 109007 597410
rect 108316 597352 108946 597408
rect 109002 597352 109007 597408
rect 108316 597350 109007 597352
rect 108316 597348 108322 597350
rect 108941 597347 109007 597350
rect 115974 597348 115980 597412
rect 116044 597410 116050 597412
rect 117221 597410 117287 597413
rect 116044 597408 117287 597410
rect 116044 597352 117226 597408
rect 117282 597352 117287 597408
rect 116044 597350 117287 597352
rect 116044 597348 116050 597350
rect 117221 597347 117287 597350
rect 120942 597348 120948 597412
rect 121012 597410 121018 597412
rect 121361 597410 121427 597413
rect 121012 597408 121427 597410
rect 121012 597352 121366 597408
rect 121422 597352 121427 597408
rect 121012 597350 121427 597352
rect 121012 597348 121018 597350
rect 121361 597347 121427 597350
rect 213545 597410 213611 597413
rect 260966 597410 260972 597412
rect 213545 597408 260972 597410
rect 213545 597352 213550 597408
rect 213606 597352 260972 597408
rect 213545 597350 260972 597352
rect 213545 597347 213611 597350
rect 260966 597348 260972 597350
rect 261036 597348 261042 597412
rect 262213 597410 262279 597413
rect 262806 597410 262812 597412
rect 262213 597408 262812 597410
rect 262213 597352 262218 597408
rect 262274 597352 262812 597408
rect 262213 597350 262812 597352
rect 262213 597347 262279 597350
rect 262806 597348 262812 597350
rect 262876 597348 262882 597412
rect 263685 597410 263751 597413
rect 263910 597410 263916 597412
rect 263685 597408 263916 597410
rect 263685 597352 263690 597408
rect 263746 597352 263916 597408
rect 263685 597350 263916 597352
rect 263685 597347 263751 597350
rect 263910 597348 263916 597350
rect 263980 597348 263986 597412
rect 266353 597410 266419 597413
rect 267590 597410 267596 597412
rect 266353 597408 267596 597410
rect 266353 597352 266358 597408
rect 266414 597352 267596 597408
rect 266353 597350 267596 597352
rect 266353 597347 266419 597350
rect 267590 597348 267596 597350
rect 267660 597348 267666 597412
rect 270401 597410 270467 597413
rect 276054 597410 276060 597412
rect 270401 597408 276060 597410
rect 270401 597352 270406 597408
rect 270462 597352 276060 597408
rect 270401 597350 276060 597352
rect 270401 597347 270467 597350
rect 276054 597348 276060 597350
rect 276124 597348 276130 597412
rect 300894 597348 300900 597412
rect 300964 597410 300970 597412
rect 357566 597410 357572 597412
rect 300964 597350 357572 597410
rect 300964 597348 300970 597350
rect 357566 597348 357572 597350
rect 357636 597348 357642 597412
rect 392669 597410 392735 597413
rect 451230 597410 451290 597486
rect 456006 597484 456012 597486
rect 456076 597484 456082 597548
rect 462313 597546 462379 597549
rect 463550 597546 463556 597548
rect 462313 597544 463556 597546
rect 462313 597488 462318 597544
rect 462374 597488 463556 597544
rect 462313 597486 463556 597488
rect 462313 597483 462379 597486
rect 463550 597484 463556 597486
rect 463620 597484 463626 597548
rect 465073 597546 465139 597549
rect 465942 597546 465948 597548
rect 465073 597544 465948 597546
rect 465073 597488 465078 597544
rect 465134 597488 465948 597544
rect 465073 597486 465948 597488
rect 465073 597483 465139 597486
rect 465942 597484 465948 597486
rect 466012 597484 466018 597548
rect 467833 597546 467899 597549
rect 468150 597546 468156 597548
rect 467833 597544 468156 597546
rect 467833 597488 467838 597544
rect 467894 597488 468156 597544
rect 467833 597486 468156 597488
rect 467833 597483 467899 597486
rect 468150 597484 468156 597486
rect 468220 597484 468226 597548
rect 473353 597546 473419 597549
rect 473486 597546 473492 597548
rect 473353 597544 473492 597546
rect 473353 597488 473358 597544
rect 473414 597488 473492 597544
rect 473353 597486 473492 597488
rect 473353 597483 473419 597486
rect 473486 597484 473492 597486
rect 473556 597484 473562 597548
rect 474733 597546 474799 597549
rect 475878 597546 475884 597548
rect 474733 597544 475884 597546
rect 474733 597488 474738 597544
rect 474794 597488 475884 597544
rect 474733 597486 475884 597488
rect 474733 597483 474799 597486
rect 475878 597484 475884 597486
rect 475948 597484 475954 597548
rect 477493 597546 477559 597549
rect 478454 597546 478460 597548
rect 477493 597544 478460 597546
rect 477493 597488 477498 597544
rect 477554 597488 478460 597544
rect 477493 597486 478460 597488
rect 477493 597483 477559 597486
rect 478454 597484 478460 597486
rect 478524 597484 478530 597548
rect 483013 597546 483079 597549
rect 483422 597546 483428 597548
rect 483013 597544 483428 597546
rect 483013 597488 483018 597544
rect 483074 597488 483428 597544
rect 483013 597486 483428 597488
rect 483013 597483 483079 597486
rect 483422 597484 483428 597486
rect 483492 597484 483498 597548
rect 485773 597546 485839 597549
rect 488533 597548 488599 597549
rect 485998 597546 486004 597548
rect 485773 597544 486004 597546
rect 485773 597488 485778 597544
rect 485834 597488 486004 597544
rect 485773 597486 486004 597488
rect 485773 597483 485839 597486
rect 485998 597484 486004 597486
rect 486068 597484 486074 597548
rect 488533 597546 488580 597548
rect 488488 597544 488580 597546
rect 488488 597488 488538 597544
rect 488488 597486 488580 597488
rect 488533 597484 488580 597486
rect 488644 597484 488650 597548
rect 495433 597546 495499 597549
rect 495934 597546 495940 597548
rect 495433 597544 495940 597546
rect 495433 597488 495438 597544
rect 495494 597488 495940 597544
rect 495433 597486 495940 597488
rect 488533 597483 488599 597484
rect 495433 597483 495499 597486
rect 495934 597484 495940 597486
rect 496004 597484 496010 597548
rect 498193 597546 498259 597549
rect 500953 597548 501019 597549
rect 498510 597546 498516 597548
rect 498193 597544 498516 597546
rect 498193 597488 498198 597544
rect 498254 597488 498516 597544
rect 498193 597486 498516 597488
rect 498193 597483 498259 597486
rect 498510 597484 498516 597486
rect 498580 597484 498586 597548
rect 500902 597484 500908 597548
rect 500972 597546 501019 597548
rect 500972 597544 501064 597546
rect 501014 597488 501064 597544
rect 500972 597486 501064 597488
rect 500972 597484 501019 597486
rect 500953 597483 501019 597484
rect 392669 597408 451290 597410
rect 392669 597352 392674 597408
rect 392730 597352 451290 597408
rect 392669 597350 451290 597352
rect 452653 597410 452719 597413
rect 453246 597410 453252 597412
rect 452653 597408 453252 597410
rect 452653 597352 452658 597408
rect 452714 597352 453252 597408
rect 452653 597350 453252 597352
rect 392669 597347 392735 597350
rect 452653 597347 452719 597350
rect 453246 597348 453252 597350
rect 453316 597348 453322 597412
rect 85573 597274 85639 597277
rect 86350 597274 86356 597276
rect 85573 597272 86356 597274
rect 85573 597216 85578 597272
rect 85634 597216 86356 597272
rect 85573 597214 86356 597216
rect 85573 597211 85639 597214
rect 86350 597212 86356 597214
rect 86420 597212 86426 597276
rect 86953 597274 87019 597277
rect 87638 597274 87644 597276
rect 86953 597272 87644 597274
rect 86953 597216 86958 597272
rect 87014 597216 87644 597272
rect 86953 597214 87644 597216
rect 86953 597211 87019 597214
rect 87638 597212 87644 597214
rect 87708 597212 87714 597276
rect 95233 597274 95299 597277
rect 95734 597274 95740 597276
rect 95233 597272 95740 597274
rect 95233 597216 95238 597272
rect 95294 597216 95740 597272
rect 95233 597214 95740 597216
rect 95233 597211 95299 597214
rect 95734 597212 95740 597214
rect 95804 597212 95810 597276
rect 99046 597274 99052 597276
rect 95926 597214 99052 597274
rect 79366 597078 84210 597138
rect 88333 597138 88399 597141
rect 88742 597138 88748 597140
rect 88333 597136 88748 597138
rect 88333 597080 88338 597136
rect 88394 597080 88748 597136
rect 88333 597078 88748 597080
rect 36997 597002 37063 597005
rect 79366 597004 79426 597078
rect 88333 597075 88399 597078
rect 88742 597076 88748 597078
rect 88812 597076 88818 597140
rect 89713 597138 89779 597141
rect 89846 597138 89852 597140
rect 89713 597136 89852 597138
rect 89713 597080 89718 597136
rect 89774 597080 89852 597136
rect 89713 597078 89852 597080
rect 89713 597075 89779 597078
rect 89846 597076 89852 597078
rect 89916 597076 89922 597140
rect 95926 597138 95986 597214
rect 99046 597212 99052 597214
rect 99116 597212 99122 597276
rect 113398 597212 113404 597276
rect 113468 597274 113474 597276
rect 114461 597274 114527 597277
rect 113468 597272 114527 597274
rect 113468 597216 114466 597272
rect 114522 597216 114527 597272
rect 113468 597214 114527 597216
rect 113468 597212 113474 597214
rect 114461 597211 114527 597214
rect 219014 597212 219020 597276
rect 219084 597274 219090 597276
rect 273478 597274 273484 597276
rect 219084 597214 273484 597274
rect 219084 597212 219090 597214
rect 273478 597212 273484 597214
rect 273548 597212 273554 597276
rect 274633 597274 274699 597277
rect 275686 597274 275692 597276
rect 274633 597272 275692 597274
rect 274633 597216 274638 597272
rect 274694 597216 275692 597272
rect 274633 597214 275692 597216
rect 274633 597211 274699 597214
rect 275686 597212 275692 597214
rect 275756 597212 275762 597276
rect 298502 597212 298508 597276
rect 298572 597274 298578 597276
rect 358854 597274 358860 597276
rect 298572 597214 358860 597274
rect 298572 597212 298578 597214
rect 358854 597212 358860 597214
rect 358924 597212 358930 597276
rect 389817 597274 389883 597277
rect 460974 597274 460980 597276
rect 389817 597272 460980 597274
rect 389817 597216 389822 597272
rect 389878 597216 460980 597272
rect 389817 597214 460980 597216
rect 389817 597211 389883 597214
rect 460974 597212 460980 597214
rect 461044 597212 461050 597276
rect 93810 597078 95986 597138
rect 96613 597138 96679 597141
rect 97022 597138 97028 597140
rect 96613 597136 97028 597138
rect 96613 597080 96618 597136
rect 96674 597080 97028 597136
rect 96613 597078 97028 597080
rect 79358 597002 79364 597004
rect 36997 597000 79364 597002
rect 36997 596944 37002 597000
rect 37058 596944 79364 597000
rect 36997 596942 79364 596944
rect 36997 596939 37063 596942
rect 79358 596940 79364 596942
rect 79428 596940 79434 597004
rect 80646 597002 80652 597004
rect 79734 596942 80652 597002
rect 36813 596866 36879 596869
rect 79734 596866 79794 596942
rect 80646 596940 80652 596942
rect 80716 597002 80722 597004
rect 93810 597002 93870 597078
rect 96613 597075 96679 597078
rect 97022 597076 97028 597078
rect 97092 597076 97098 597140
rect 125910 597076 125916 597140
rect 125980 597138 125986 597140
rect 126881 597138 126947 597141
rect 125980 597136 126947 597138
rect 125980 597080 126886 597136
rect 126942 597080 126947 597136
rect 125980 597078 126947 597080
rect 125980 597076 125986 597078
rect 126881 597075 126947 597078
rect 138422 597076 138428 597140
rect 138492 597138 138498 597140
rect 139301 597138 139367 597141
rect 138492 597136 139367 597138
rect 138492 597080 139306 597136
rect 139362 597080 139367 597136
rect 138492 597078 139367 597080
rect 138492 597076 138498 597078
rect 139301 597075 139367 597078
rect 219985 597138 220051 597141
rect 270401 597138 270467 597141
rect 219985 597136 270467 597138
rect 219985 597080 219990 597136
rect 220046 597080 270406 597136
rect 270462 597080 270467 597136
rect 219985 597078 270467 597080
rect 219985 597075 220051 597078
rect 270401 597075 270467 597078
rect 270585 597138 270651 597141
rect 273253 597140 273319 597141
rect 271086 597138 271092 597140
rect 270585 597136 271092 597138
rect 270585 597080 270590 597136
rect 270646 597080 271092 597136
rect 270585 597078 271092 597080
rect 270585 597075 270651 597078
rect 271086 597076 271092 597078
rect 271156 597076 271162 597140
rect 273253 597138 273300 597140
rect 273208 597136 273300 597138
rect 273208 597080 273258 597136
rect 273208 597078 273300 597080
rect 273253 597076 273300 597078
rect 273364 597076 273370 597140
rect 287053 597138 287119 597141
rect 288198 597138 288204 597140
rect 287053 597136 288204 597138
rect 287053 597080 287058 597136
rect 287114 597080 288204 597136
rect 287053 597078 288204 597080
rect 273253 597075 273319 597076
rect 287053 597075 287119 597078
rect 288198 597076 288204 597078
rect 288268 597076 288274 597140
rect 357014 597076 357020 597140
rect 357084 597138 357090 597140
rect 438526 597138 438532 597140
rect 357084 597078 438532 597138
rect 357084 597076 357090 597078
rect 438526 597076 438532 597078
rect 438596 597076 438602 597140
rect 440325 597138 440391 597141
rect 440734 597138 440740 597140
rect 440325 597136 440740 597138
rect 440325 597080 440330 597136
rect 440386 597080 440740 597136
rect 440325 597078 440740 597080
rect 440325 597075 440391 597078
rect 440734 597076 440740 597078
rect 440804 597138 440810 597140
rect 459134 597138 459140 597140
rect 440804 597078 459140 597138
rect 440804 597076 440810 597078
rect 459134 597076 459140 597078
rect 459204 597076 459210 597140
rect 80716 596942 93870 597002
rect 80716 596940 80722 596942
rect 111006 596940 111012 597004
rect 111076 597002 111082 597004
rect 111701 597002 111767 597005
rect 118601 597004 118667 597005
rect 111076 597000 111767 597002
rect 111076 596944 111706 597000
rect 111762 596944 111767 597000
rect 111076 596942 111767 596944
rect 111076 596940 111082 596942
rect 111701 596939 111767 596942
rect 118550 596940 118556 597004
rect 118620 597002 118667 597004
rect 118620 597000 118712 597002
rect 118662 596944 118712 597000
rect 118620 596942 118712 596944
rect 118620 596940 118667 596942
rect 141918 596940 141924 597004
rect 141988 597002 141994 597004
rect 177205 597002 177271 597005
rect 141988 597000 177271 597002
rect 141988 596944 177210 597000
rect 177266 596944 177271 597000
rect 141988 596942 177271 596944
rect 141988 596940 141994 596942
rect 118601 596939 118667 596940
rect 177205 596939 177271 596942
rect 211061 597002 211127 597005
rect 277301 597002 277367 597005
rect 211061 597000 277367 597002
rect 211061 596944 211066 597000
rect 211122 596944 277306 597000
rect 277362 596944 277367 597000
rect 211061 596942 277367 596944
rect 211061 596939 211127 596942
rect 277301 596939 277367 596942
rect 325918 596940 325924 597004
rect 325988 597002 325994 597004
rect 326981 597002 327047 597005
rect 441613 597004 441679 597005
rect 325988 597000 327047 597002
rect 325988 596944 326986 597000
rect 327042 596944 327047 597000
rect 325988 596942 327047 596944
rect 325988 596940 325994 596942
rect 326981 596939 327047 596942
rect 356646 596940 356652 597004
rect 356716 597002 356722 597004
rect 441102 597002 441108 597004
rect 356716 596942 441108 597002
rect 356716 596940 356722 596942
rect 441102 596940 441108 596942
rect 441172 596940 441178 597004
rect 441613 597000 441660 597004
rect 441724 597002 441730 597004
rect 445845 597002 445911 597005
rect 446254 597002 446260 597004
rect 441613 596944 441618 597000
rect 441613 596940 441660 596944
rect 441724 596942 441770 597002
rect 445845 597000 446260 597002
rect 445845 596944 445850 597000
rect 445906 596944 446260 597000
rect 445845 596942 446260 596944
rect 441724 596940 441730 596942
rect 441613 596939 441679 596940
rect 445845 596939 445911 596942
rect 446254 596940 446260 596942
rect 446324 596940 446330 597004
rect 447225 597002 447291 597005
rect 447542 597002 447548 597004
rect 447225 597000 447548 597002
rect 447225 596944 447230 597000
rect 447286 596944 447548 597000
rect 447225 596942 447548 596944
rect 447225 596939 447291 596942
rect 447542 596940 447548 596942
rect 447612 596940 447618 597004
rect 448513 597002 448579 597005
rect 448646 597002 448652 597004
rect 448513 597000 448652 597002
rect 448513 596944 448518 597000
rect 448574 596944 448652 597000
rect 448513 596942 448652 596944
rect 448513 596939 448579 596942
rect 448646 596940 448652 596942
rect 448716 596940 448722 597004
rect 454033 597002 454099 597005
rect 454350 597002 454356 597004
rect 454033 597000 454356 597002
rect 454033 596944 454038 597000
rect 454094 596944 454356 597000
rect 454033 596942 454356 596944
rect 454033 596939 454099 596942
rect 454350 596940 454356 596942
rect 454420 596940 454426 597004
rect 455413 597002 455479 597005
rect 455638 597002 455644 597004
rect 455413 597000 455644 597002
rect 455413 596944 455418 597000
rect 455474 596944 455644 597000
rect 455413 596942 455644 596944
rect 455413 596939 455479 596942
rect 455638 596940 455644 596942
rect 455708 596940 455714 597004
rect 480253 597002 480319 597005
rect 480846 597002 480852 597004
rect 480253 597000 480852 597002
rect 480253 596944 480258 597000
rect 480314 596944 480852 597000
rect 480253 596942 480852 596944
rect 480253 596939 480319 596942
rect 480846 596940 480852 596942
rect 480916 596940 480922 597004
rect 502333 597002 502399 597005
rect 503294 597002 503300 597004
rect 502333 597000 503300 597002
rect 502333 596944 502338 597000
rect 502394 596944 503300 597000
rect 502333 596942 503300 596944
rect 502333 596939 502399 596942
rect 503294 596940 503300 596942
rect 503364 596940 503370 597004
rect 82813 596868 82879 596869
rect 82813 596866 82860 596868
rect 36813 596864 79794 596866
rect 36813 596808 36818 596864
rect 36874 596808 79794 596864
rect 36813 596806 79794 596808
rect 82768 596864 82860 596866
rect 82768 596808 82818 596864
rect 82768 596806 82860 596808
rect 36813 596803 36879 596806
rect 82813 596804 82860 596806
rect 82924 596804 82930 596868
rect 103278 596804 103284 596868
rect 103348 596866 103354 596868
rect 219934 596866 219940 596868
rect 103348 596806 219940 596866
rect 103348 596804 103354 596806
rect 219934 596804 219940 596806
rect 220004 596804 220010 596868
rect 238518 596804 238524 596868
rect 238588 596866 238594 596868
rect 238753 596866 238819 596869
rect 238588 596864 238819 596866
rect 238588 596808 238758 596864
rect 238814 596808 238819 596864
rect 238588 596806 238819 596808
rect 238588 596804 238594 596806
rect 82813 596803 82879 596804
rect 238753 596803 238819 596806
rect 240133 596866 240199 596869
rect 240542 596866 240548 596868
rect 240133 596864 240548 596866
rect 240133 596808 240138 596864
rect 240194 596808 240548 596864
rect 240133 596806 240548 596808
rect 240133 596803 240199 596806
rect 240542 596804 240548 596806
rect 240612 596804 240618 596868
rect 241513 596866 241579 596869
rect 241646 596866 241652 596868
rect 241513 596864 241652 596866
rect 241513 596808 241518 596864
rect 241574 596808 241652 596864
rect 241513 596806 241652 596808
rect 241513 596803 241579 596806
rect 241646 596804 241652 596806
rect 241716 596804 241722 596868
rect 247125 596866 247191 596869
rect 247534 596866 247540 596868
rect 247125 596864 247540 596866
rect 247125 596808 247130 596864
rect 247186 596808 247540 596864
rect 247125 596806 247540 596808
rect 247125 596803 247191 596806
rect 247534 596804 247540 596806
rect 247604 596804 247610 596868
rect 249885 596866 249951 596869
rect 250110 596866 250116 596868
rect 249885 596864 250116 596866
rect 249885 596808 249890 596864
rect 249946 596808 250116 596864
rect 249885 596806 250116 596808
rect 249885 596803 249951 596806
rect 250110 596804 250116 596806
rect 250180 596804 250186 596868
rect 251398 596804 251404 596868
rect 251468 596866 251474 596868
rect 252185 596866 252251 596869
rect 251468 596864 252251 596866
rect 251468 596808 252190 596864
rect 252246 596808 252251 596864
rect 251468 596806 252251 596808
rect 251468 596804 251474 596806
rect 252185 596803 252251 596806
rect 265065 596866 265131 596869
rect 265198 596866 265204 596868
rect 265065 596864 265204 596866
rect 265065 596808 265070 596864
rect 265126 596808 265204 596864
rect 265065 596806 265204 596808
rect 265065 596803 265131 596806
rect 265198 596804 265204 596806
rect 265268 596804 265274 596868
rect 278078 596866 278084 596868
rect 267690 596806 278084 596866
rect 55397 596730 55463 596733
rect 55990 596730 55996 596732
rect 55397 596728 55996 596730
rect 55397 596672 55402 596728
rect 55458 596672 55996 596728
rect 55397 596670 55996 596672
rect 55397 596667 55463 596670
rect 55990 596668 55996 596670
rect 56060 596668 56066 596732
rect 100886 596668 100892 596732
rect 100956 596730 100962 596732
rect 102041 596730 102107 596733
rect 100956 596728 102107 596730
rect 100956 596672 102046 596728
rect 102102 596672 102107 596728
rect 100956 596670 102107 596672
rect 100956 596668 100962 596670
rect 102041 596667 102107 596670
rect 216581 596730 216647 596733
rect 259545 596732 259611 596733
rect 257838 596730 257844 596732
rect 216581 596728 257844 596730
rect 216581 596672 216586 596728
rect 216642 596672 257844 596728
rect 216581 596670 257844 596672
rect 216581 596667 216647 596670
rect 257838 596668 257844 596670
rect 257908 596668 257914 596732
rect 259494 596730 259500 596732
rect 259418 596670 259500 596730
rect 259564 596730 259611 596732
rect 267690 596730 267750 596806
rect 278078 596804 278084 596806
rect 278148 596804 278154 596868
rect 311014 596804 311020 596868
rect 311084 596866 311090 596868
rect 311801 596866 311867 596869
rect 311084 596864 311867 596866
rect 311084 596808 311806 596864
rect 311862 596808 311867 596864
rect 311084 596806 311867 596808
rect 311084 596804 311090 596806
rect 311801 596803 311867 596806
rect 320950 596804 320956 596868
rect 321020 596866 321026 596868
rect 321461 596866 321527 596869
rect 321020 596864 321527 596866
rect 321020 596808 321466 596864
rect 321522 596808 321527 596864
rect 321020 596806 321527 596808
rect 321020 596804 321026 596806
rect 321461 596803 321527 596806
rect 323342 596804 323348 596868
rect 323412 596866 323418 596868
rect 324221 596866 324287 596869
rect 323412 596864 324287 596866
rect 323412 596808 324226 596864
rect 324282 596808 324287 596864
rect 323412 596806 324287 596808
rect 323412 596804 323418 596806
rect 324221 596803 324287 596806
rect 356789 596866 356855 596869
rect 458398 596866 458404 596868
rect 356789 596864 458404 596866
rect 356789 596808 356794 596864
rect 356850 596808 458404 596864
rect 356789 596806 458404 596808
rect 356789 596803 356855 596806
rect 458398 596804 458404 596806
rect 458468 596804 458474 596868
rect 505093 596866 505159 596869
rect 505870 596866 505876 596868
rect 505093 596864 505876 596866
rect 505093 596808 505098 596864
rect 505154 596808 505876 596864
rect 505093 596806 505876 596808
rect 505093 596803 505159 596806
rect 505870 596804 505876 596806
rect 505940 596804 505946 596868
rect 259564 596728 267750 596730
rect 259606 596672 267750 596728
rect 259494 596668 259500 596670
rect 259564 596670 267750 596672
rect 267917 596730 267983 596733
rect 268694 596730 268700 596732
rect 267917 596728 268700 596730
rect 267917 596672 267922 596728
rect 267978 596672 268700 596728
rect 267917 596670 268700 596672
rect 259564 596668 259611 596670
rect 259545 596667 259611 596668
rect 267917 596667 267983 596670
rect 268694 596668 268700 596670
rect 268764 596668 268770 596732
rect 269113 596730 269179 596733
rect 269798 596730 269804 596732
rect 269113 596728 269804 596730
rect 269113 596672 269118 596728
rect 269174 596672 269804 596728
rect 269113 596670 269804 596672
rect 269113 596667 269179 596670
rect 269798 596668 269804 596670
rect 269868 596668 269874 596732
rect 313406 596668 313412 596732
rect 313476 596730 313482 596732
rect 314561 596730 314627 596733
rect 313476 596728 314627 596730
rect 313476 596672 314566 596728
rect 314622 596672 314627 596728
rect 313476 596670 314627 596672
rect 313476 596668 313482 596670
rect 314561 596667 314627 596670
rect 318558 596668 318564 596732
rect 318628 596730 318634 596732
rect 318701 596730 318767 596733
rect 419533 596732 419599 596733
rect 419533 596730 419580 596732
rect 318628 596728 318767 596730
rect 318628 596672 318706 596728
rect 318762 596672 318767 596728
rect 318628 596670 318767 596672
rect 419488 596728 419580 596730
rect 419488 596672 419538 596728
rect 419488 596670 419580 596672
rect 318628 596668 318634 596670
rect 318701 596667 318767 596670
rect 419533 596668 419580 596670
rect 419644 596668 419650 596732
rect 427813 596730 427879 596733
rect 428222 596730 428228 596732
rect 427813 596728 428228 596730
rect 427813 596672 427818 596728
rect 427874 596672 428228 596728
rect 427813 596670 428228 596672
rect 419533 596667 419599 596668
rect 427813 596667 427879 596670
rect 428222 596668 428228 596670
rect 428292 596668 428298 596732
rect 430665 596730 430731 596733
rect 431953 596732 432019 596733
rect 433425 596732 433491 596733
rect 431166 596730 431172 596732
rect 430665 596728 431172 596730
rect 430665 596672 430670 596728
rect 430726 596672 431172 596728
rect 430665 596670 431172 596672
rect 430665 596667 430731 596670
rect 431166 596668 431172 596670
rect 431236 596668 431242 596732
rect 431902 596668 431908 596732
rect 431972 596730 432019 596732
rect 433374 596730 433380 596732
rect 431972 596728 432064 596730
rect 432014 596672 432064 596728
rect 431972 596670 432064 596672
rect 433334 596670 433380 596730
rect 433444 596728 433491 596732
rect 433486 596672 433491 596728
rect 431972 596668 432019 596670
rect 433374 596668 433380 596670
rect 433444 596668 433491 596672
rect 431953 596667 432019 596668
rect 433425 596667 433491 596668
rect 438853 596730 438919 596733
rect 458030 596730 458036 596732
rect 438853 596728 458036 596730
rect 438853 596672 438858 596728
rect 438914 596672 458036 596728
rect 438853 596670 458036 596672
rect 438853 596667 438919 596670
rect 458030 596668 458036 596670
rect 458100 596668 458106 596732
rect 492673 596730 492739 596733
rect 493358 596730 493364 596732
rect 492673 596728 493364 596730
rect 492673 596672 492678 596728
rect 492734 596672 493364 596728
rect 492673 596670 493364 596672
rect 492673 596667 492739 596670
rect 493358 596668 493364 596670
rect 493428 596668 493434 596732
rect 91185 596594 91251 596597
rect 92238 596594 92244 596596
rect 91185 596592 92244 596594
rect 91185 596536 91190 596592
rect 91246 596536 92244 596592
rect 91185 596534 92244 596536
rect 91185 596531 91251 596534
rect 92238 596532 92244 596534
rect 92308 596532 92314 596596
rect 94037 596594 94103 596597
rect 94446 596594 94452 596596
rect 94037 596592 94452 596594
rect 94037 596536 94042 596592
rect 94098 596536 94452 596592
rect 94037 596534 94452 596536
rect 94037 596531 94103 596534
rect 94446 596532 94452 596534
rect 94516 596532 94522 596596
rect 106038 596532 106044 596596
rect 106108 596594 106114 596596
rect 106181 596594 106247 596597
rect 106108 596592 106247 596594
rect 106108 596536 106186 596592
rect 106242 596536 106247 596592
rect 106108 596534 106247 596536
rect 106108 596532 106114 596534
rect 106181 596531 106247 596534
rect 216254 596532 216260 596596
rect 216324 596594 216330 596596
rect 255998 596594 256004 596596
rect 216324 596534 256004 596594
rect 216324 596532 216330 596534
rect 255998 596532 256004 596534
rect 256068 596532 256074 596596
rect 259453 596594 259519 596597
rect 260598 596594 260604 596596
rect 259453 596592 260604 596594
rect 259453 596536 259458 596592
rect 259514 596536 260604 596592
rect 259453 596534 260604 596536
rect 259453 596531 259519 596534
rect 260598 596532 260604 596534
rect 260668 596594 260674 596596
rect 279182 596594 279188 596596
rect 260668 596534 279188 596594
rect 260668 596532 260674 596534
rect 279182 596532 279188 596534
rect 279252 596532 279258 596596
rect 315798 596532 315804 596596
rect 315868 596594 315874 596596
rect 315941 596594 316007 596597
rect 453614 596594 453620 596596
rect 315868 596592 316007 596594
rect 315868 596536 315946 596592
rect 316002 596536 316007 596592
rect 315868 596534 316007 596536
rect 315868 596532 315874 596534
rect 315941 596531 316007 596534
rect 446384 596534 453620 596594
rect 83590 596396 83596 596460
rect 83660 596458 83666 596460
rect 84101 596458 84167 596461
rect 91093 596460 91159 596461
rect 91093 596458 91140 596460
rect 83660 596456 84167 596458
rect 83660 596400 84106 596456
rect 84162 596400 84167 596456
rect 83660 596398 84167 596400
rect 91048 596456 91140 596458
rect 91048 596400 91098 596456
rect 91048 596398 91140 596400
rect 83660 596396 83666 596398
rect 84101 596395 84167 596398
rect 91093 596396 91140 596398
rect 91204 596396 91210 596460
rect 96102 596396 96108 596460
rect 96172 596458 96178 596460
rect 96521 596458 96587 596461
rect 96172 596456 96587 596458
rect 96172 596400 96526 596456
rect 96582 596400 96587 596456
rect 96172 596398 96587 596400
rect 96172 596396 96178 596398
rect 91093 596395 91159 596396
rect 96521 596395 96587 596398
rect 98494 596396 98500 596460
rect 98564 596458 98570 596460
rect 99281 596458 99347 596461
rect 266353 596460 266419 596461
rect 98564 596456 99347 596458
rect 98564 596400 99286 596456
rect 99342 596400 99347 596456
rect 98564 596398 99347 596400
rect 98564 596396 98570 596398
rect 99281 596395 99347 596398
rect 266302 596396 266308 596460
rect 266372 596458 266419 596460
rect 271873 596458 271939 596461
rect 306097 596460 306163 596461
rect 272190 596458 272196 596460
rect 266372 596456 266464 596458
rect 266414 596400 266464 596456
rect 266372 596398 266464 596400
rect 271873 596456 272196 596458
rect 271873 596400 271878 596456
rect 271934 596400 272196 596456
rect 271873 596398 272196 596400
rect 266372 596396 266419 596398
rect 266353 596395 266419 596396
rect 271873 596395 271939 596398
rect 272190 596396 272196 596398
rect 272260 596396 272266 596460
rect 306046 596396 306052 596460
rect 306116 596458 306163 596460
rect 306116 596456 306208 596458
rect 306158 596400 306208 596456
rect 306116 596398 306208 596400
rect 306116 596396 306163 596398
rect 308622 596396 308628 596460
rect 308692 596458 308698 596460
rect 309041 596458 309107 596461
rect 308692 596456 309107 596458
rect 308692 596400 309046 596456
rect 309102 596400 309107 596456
rect 308692 596398 309107 596400
rect 308692 596396 308698 596398
rect 306097 596395 306163 596396
rect 309041 596395 309107 596398
rect 392853 596458 392919 596461
rect 446384 596458 446444 596534
rect 453614 596532 453620 596534
rect 453684 596532 453690 596596
rect 392853 596456 446444 596458
rect 392853 596400 392858 596456
rect 392914 596400 446444 596456
rect 392853 596398 446444 596400
rect 449985 596458 450051 596461
rect 450854 596458 450860 596460
rect 449985 596456 450860 596458
rect 449985 596400 449990 596456
rect 450046 596400 450860 596456
rect 449985 596398 450860 596400
rect 392853 596395 392919 596398
rect 449985 596395 450051 596398
rect 450854 596396 450860 596398
rect 450924 596396 450930 596460
rect 451089 596458 451155 596461
rect 451273 596458 451339 596461
rect 451089 596456 451339 596458
rect 451089 596400 451094 596456
rect 451150 596400 451278 596456
rect 451334 596400 451339 596456
rect 451089 596398 451339 596400
rect 451089 596395 451155 596398
rect 451273 596395 451339 596398
rect 91001 596324 91067 596325
rect 90950 596260 90956 596324
rect 91020 596322 91067 596324
rect 91020 596320 91112 596322
rect 91062 596264 91112 596320
rect 91020 596262 91112 596264
rect 91020 596260 91067 596262
rect 210734 596260 210740 596324
rect 210804 596322 210810 596324
rect 253606 596322 253612 596324
rect 210804 596262 253612 596322
rect 210804 596260 210810 596262
rect 253606 596260 253612 596262
rect 253676 596260 253682 596324
rect 273253 596322 273319 596325
rect 274398 596322 274404 596324
rect 273253 596320 274404 596322
rect 273253 596264 273258 596320
rect 273314 596264 274404 596320
rect 273253 596262 274404 596264
rect 91001 596259 91067 596260
rect 273253 596259 273319 596262
rect 274398 596260 274404 596262
rect 274468 596260 274474 596324
rect 295926 596260 295932 596324
rect 295996 596322 296002 596324
rect 296345 596322 296411 596325
rect 303521 596324 303587 596325
rect 295996 596320 296411 596322
rect 295996 596264 296350 596320
rect 296406 596264 296411 596320
rect 295996 596262 296411 596264
rect 295996 596260 296002 596262
rect 296345 596259 296411 596262
rect 303470 596260 303476 596324
rect 303540 596322 303587 596324
rect 448513 596322 448579 596325
rect 449750 596322 449756 596324
rect 303540 596320 303632 596322
rect 303582 596264 303632 596320
rect 303540 596262 303632 596264
rect 448513 596320 449756 596322
rect 448513 596264 448518 596320
rect 448574 596264 449756 596320
rect 448513 596262 449756 596264
rect 303540 596260 303587 596262
rect 303521 596259 303587 596260
rect 448513 596259 448579 596262
rect 449750 596260 449756 596262
rect 449820 596260 449826 596324
rect 456793 596322 456859 596325
rect 456926 596322 456932 596324
rect 456793 596320 456932 596322
rect 456793 596264 456798 596320
rect 456854 596264 456932 596320
rect 456793 596262 456932 596264
rect 456793 596259 456859 596262
rect 456926 596260 456932 596262
rect 456996 596260 457002 596324
rect 470358 596260 470364 596324
rect 470428 596322 470434 596324
rect 470593 596322 470659 596325
rect 470428 596320 470659 596322
rect 470428 596264 470598 596320
rect 470654 596264 470659 596320
rect 470428 596262 470659 596264
rect 470428 596260 470434 596262
rect 470593 596259 470659 596262
rect 489678 596260 489684 596324
rect 489748 596322 489754 596324
rect 489913 596322 489979 596325
rect 489748 596320 489979 596322
rect 489748 596264 489918 596320
rect 489974 596264 489979 596320
rect 489748 596262 489979 596264
rect 489748 596260 489754 596262
rect 489913 596259 489979 596262
rect 213637 594554 213703 594557
rect 263593 594554 263659 594557
rect 213637 594552 263659 594554
rect 213637 594496 213642 594552
rect 213698 594496 263598 594552
rect 263654 594496 263659 594552
rect 213637 594494 263659 594496
rect 213637 594491 213703 594494
rect 263593 594491 263659 594494
rect 399334 594492 399340 594556
rect 399404 594554 399410 594556
rect 442993 594554 443059 594557
rect 399404 594552 443059 594554
rect 399404 594496 442998 594552
rect 443054 594496 443059 594552
rect 399404 594494 443059 594496
rect 399404 594492 399410 594494
rect 442993 594491 443059 594494
rect 213729 594418 213795 594421
rect 264973 594418 265039 594421
rect 213729 594416 265039 594418
rect 213729 594360 213734 594416
rect 213790 594360 264978 594416
rect 265034 594360 265039 594416
rect 213729 594358 265039 594360
rect 213729 594355 213795 594358
rect 264973 594355 265039 594358
rect 390093 594418 390159 594421
rect 462313 594418 462379 594421
rect 390093 594416 462379 594418
rect 390093 594360 390098 594416
rect 390154 594360 462318 594416
rect 462374 594360 462379 594416
rect 390093 594358 462379 594360
rect 390093 594355 390159 594358
rect 462313 594355 462379 594358
rect 213821 594282 213887 594285
rect 267733 594282 267799 594285
rect 213821 594280 267799 594282
rect 213821 594224 213826 594280
rect 213882 594224 267738 594280
rect 267794 594224 267799 594280
rect 213821 594222 267799 594224
rect 213821 594219 213887 594222
rect 267733 594219 267799 594222
rect 390461 594282 390527 594285
rect 465073 594282 465139 594285
rect 390461 594280 465139 594282
rect 390461 594224 390466 594280
rect 390522 594224 465078 594280
rect 465134 594224 465139 594280
rect 390461 594222 465139 594224
rect 390461 594219 390527 594222
rect 465073 594219 465139 594222
rect 215150 594084 215156 594148
rect 215220 594146 215226 594148
rect 270493 594146 270559 594149
rect 215220 594144 270559 594146
rect 215220 594088 270498 594144
rect 270554 594088 270559 594144
rect 215220 594086 270559 594088
rect 215220 594084 215226 594086
rect 270493 594083 270559 594086
rect 390277 594146 390343 594149
rect 467833 594146 467899 594149
rect 390277 594144 467899 594146
rect 390277 594088 390282 594144
rect 390338 594088 467838 594144
rect 467894 594088 467899 594144
rect 390277 594086 467899 594088
rect 390277 594083 390343 594086
rect 467833 594083 467899 594086
rect 217726 593948 217732 594012
rect 217796 594010 217802 594012
rect 282913 594010 282979 594013
rect 217796 594008 282979 594010
rect 217796 593952 282918 594008
rect 282974 593952 282979 594008
rect 217796 593950 282979 593952
rect 217796 593948 217802 593950
rect 282913 593947 282979 593950
rect 389725 594010 389791 594013
rect 470593 594010 470659 594013
rect 389725 594008 470659 594010
rect 389725 593952 389730 594008
rect 389786 593952 470598 594008
rect 470654 593952 470659 594008
rect 389725 593950 470659 593952
rect 389725 593947 389791 593950
rect 470593 593947 470659 593950
rect -960 592908 480 593148
rect 358118 592588 358124 592652
rect 358188 592650 358194 592652
rect 505093 592650 505159 592653
rect 358188 592648 505159 592650
rect 358188 592592 505098 592648
rect 505154 592592 505159 592648
rect 358188 592590 505159 592592
rect 358188 592588 358194 592590
rect 505093 592587 505159 592590
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 2773 580002 2839 580005
rect -960 580000 2839 580002
rect -960 579944 2778 580000
rect 2834 579944 2839 580000
rect -960 579942 2839 579944
rect -960 579852 480 579942
rect 2773 579939 2839 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect 212390 571916 212396 571980
rect 212460 571978 212466 571980
rect 427813 571978 427879 571981
rect 212460 571976 427879 571978
rect 212460 571920 427818 571976
rect 427874 571920 427879 571976
rect 212460 571918 427879 571920
rect 212460 571916 212466 571918
rect 427813 571915 427879 571918
rect 74441 570754 74507 570757
rect 218646 570754 218652 570756
rect 74441 570752 218652 570754
rect 74441 570696 74446 570752
rect 74502 570696 218652 570752
rect 74441 570694 218652 570696
rect 74441 570691 74507 570694
rect 218646 570692 218652 570694
rect 218716 570692 218722 570756
rect 216438 570556 216444 570620
rect 216508 570618 216514 570620
rect 430573 570618 430639 570621
rect 216508 570616 430639 570618
rect 216508 570560 430578 570616
rect 430634 570560 430639 570616
rect 216508 570558 430639 570560
rect 216508 570556 216514 570558
rect 430573 570555 430639 570558
rect 213913 567218 213979 567221
rect 217910 567218 217916 567220
rect 213913 567216 217916 567218
rect 213913 567160 213918 567216
rect 213974 567160 217916 567216
rect 213913 567158 217916 567160
rect 213913 567155 213979 567158
rect 217910 567156 217916 567158
rect 217980 567156 217986 567220
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 210918 566476 210924 566540
rect 210988 566538 210994 566540
rect 247033 566538 247099 566541
rect 210988 566536 247099 566538
rect 210988 566480 247038 566536
rect 247094 566480 247099 566536
rect 210988 566478 247099 566480
rect 210988 566476 210994 566478
rect 247033 566475 247099 566478
rect 71681 566402 71747 566405
rect 212574 566402 212580 566404
rect 71681 566400 212580 566402
rect 71681 566344 71686 566400
rect 71742 566344 212580 566400
rect 71681 566342 212580 566344
rect 71681 566339 71747 566342
rect 212574 566340 212580 566342
rect 212644 566340 212650 566404
rect 170857 565860 170923 565861
rect 170806 565858 170812 565860
rect 170766 565798 170812 565858
rect 170876 565856 170923 565860
rect 170918 565800 170923 565856
rect 170806 565796 170812 565798
rect 170876 565796 170923 565800
rect 350942 565796 350948 565860
rect 351012 565858 351018 565860
rect 351085 565858 351151 565861
rect 530945 565860 531011 565861
rect 530894 565858 530900 565860
rect 351012 565856 351151 565858
rect 351012 565800 351090 565856
rect 351146 565800 351151 565856
rect 351012 565798 351151 565800
rect 530854 565798 530900 565858
rect 530964 565856 531011 565860
rect 531006 565800 531011 565856
rect 351012 565796 351018 565798
rect 170857 565795 170923 565796
rect 351085 565795 351151 565798
rect 530894 565796 530900 565798
rect 530964 565796 531011 565800
rect 530945 565795 531011 565796
rect 146201 565450 146267 565453
rect 203374 565450 203380 565452
rect 146201 565448 203380 565450
rect 146201 565392 146206 565448
rect 146262 565392 203380 565448
rect 146201 565390 203380 565392
rect 146201 565387 146267 565390
rect 203374 565388 203380 565390
rect 203444 565388 203450 565452
rect 129641 565314 129707 565317
rect 206134 565314 206140 565316
rect 129641 565312 206140 565314
rect 129641 565256 129646 565312
rect 129702 565256 206140 565312
rect 129641 565254 206140 565256
rect 129641 565251 129707 565254
rect 206134 565252 206140 565254
rect 206204 565252 206210 565316
rect 93761 565178 93827 565181
rect 206318 565178 206324 565180
rect 93761 565176 206324 565178
rect 93761 565120 93766 565176
rect 93822 565120 206324 565176
rect 93761 565118 206324 565120
rect 93761 565115 93827 565118
rect 206318 565116 206324 565118
rect 206388 565116 206394 565180
rect 68921 565042 68987 565045
rect 208710 565042 208716 565044
rect 68921 565040 208716 565042
rect 68921 564984 68926 565040
rect 68982 564984 208716 565040
rect 68921 564982 208716 564984
rect 68921 564979 68987 564982
rect 208710 564980 208716 564982
rect 208780 564980 208786 565044
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect 219750 563620 219756 563684
rect 219820 563682 219826 563684
rect 433333 563682 433399 563685
rect 219820 563680 433399 563682
rect 219820 563624 433338 563680
rect 433394 563624 433399 563680
rect 219820 563622 433399 563624
rect 219820 563620 219826 563622
rect 433333 563619 433399 563622
rect 178493 560282 178559 560285
rect 179045 560282 179111 560285
rect 178493 560280 179111 560282
rect 178493 560224 178498 560280
rect 178554 560224 179050 560280
rect 179106 560224 179111 560280
rect 178493 560222 179111 560224
rect 178493 560219 178559 560222
rect 179045 560219 179111 560222
rect 358813 560282 358879 560285
rect 359733 560282 359799 560285
rect 358813 560280 359799 560282
rect 358813 560224 358818 560280
rect 358874 560224 359738 560280
rect 359794 560224 359799 560280
rect 358813 560222 359799 560224
rect 358813 560219 358879 560222
rect 359733 560219 359799 560222
rect 176548 559194 177130 559220
rect 179045 559194 179111 559197
rect 359733 559194 359799 559197
rect 538213 559194 538279 559197
rect 176548 559192 179111 559194
rect 176548 559160 179050 559192
rect 177070 559136 179050 559160
rect 179106 559136 179111 559192
rect 177070 559134 179111 559136
rect 356562 559192 359799 559194
rect 356562 559136 359738 559192
rect 359794 559136 359799 559192
rect 356562 559134 359799 559136
rect 536558 559192 538279 559194
rect 536558 559136 538218 559192
rect 538274 559136 538279 559192
rect 536558 559134 538279 559136
rect 179045 559131 179111 559134
rect 359733 559131 359799 559134
rect 538213 559131 538279 559134
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 37825 517442 37891 517445
rect 37825 517440 40050 517442
rect 37825 517384 37830 517440
rect 37886 517384 40050 517440
rect 37825 517382 40050 517384
rect 37825 517379 37891 517382
rect 39990 516894 40050 517382
rect 217225 516898 217291 516901
rect 219390 516898 220064 516924
rect 217225 516896 220064 516898
rect 217225 516840 217230 516896
rect 217286 516864 220064 516896
rect 397269 516898 397335 516901
rect 399342 516898 400016 516924
rect 397269 516896 400016 516898
rect 217286 516840 219450 516864
rect 217225 516838 219450 516840
rect 397269 516840 397274 516896
rect 397330 516864 400016 516896
rect 397330 516840 399402 516864
rect 397269 516838 399402 516840
rect 217225 516835 217291 516838
rect 397269 516835 397335 516838
rect 216765 516218 216831 516221
rect 217225 516218 217291 516221
rect 216765 516216 217291 516218
rect 216765 516160 216770 516216
rect 216826 516160 217230 516216
rect 217286 516160 217291 516216
rect 216765 516158 217291 516160
rect 216765 516155 216831 516158
rect 217225 516155 217291 516158
rect 396441 516218 396507 516221
rect 397269 516218 397335 516221
rect 396441 516216 397335 516218
rect 396441 516160 396446 516216
rect 396502 516160 397274 516216
rect 397330 516160 397335 516216
rect 396441 516158 397335 516160
rect 396441 516155 396507 516158
rect 397269 516155 397335 516158
rect 37733 516082 37799 516085
rect 37733 516080 40050 516082
rect 37733 516024 37738 516080
rect 37794 516024 40050 516080
rect 37733 516022 40050 516024
rect 37733 516019 37799 516022
rect 39990 515942 40050 516022
rect 216949 515946 217015 515949
rect 217133 515946 217199 515949
rect 219390 515946 220064 515972
rect 216949 515944 220064 515946
rect 216949 515888 216954 515944
rect 217010 515888 217138 515944
rect 217194 515912 220064 515944
rect 396901 515946 396967 515949
rect 399342 515946 400016 515972
rect 396901 515944 400016 515946
rect 217194 515888 219450 515912
rect 216949 515886 219450 515888
rect 396901 515888 396906 515944
rect 396962 515912 400016 515944
rect 396962 515888 399402 515912
rect 396901 515886 399402 515888
rect 216949 515883 217015 515886
rect 217133 515883 217199 515886
rect 396901 515883 396967 515886
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 396533 514858 396599 514861
rect 396901 514858 396967 514861
rect 396533 514856 396967 514858
rect 396533 514800 396538 514856
rect 396594 514800 396906 514856
rect 396962 514800 396967 514856
rect 396533 514798 396967 514800
rect 396533 514795 396599 514798
rect 396901 514795 396967 514798
rect 38469 514044 38535 514045
rect 38469 514042 38516 514044
rect 38388 514040 38516 514042
rect 38580 514042 38586 514044
rect 38388 513984 38474 514040
rect 38388 513982 38516 513984
rect 38469 513980 38516 513982
rect 38580 513982 40050 514042
rect 38580 513980 38586 513982
rect 38469 513979 38535 513980
rect 39990 513766 40050 513982
rect 217041 513770 217107 513773
rect 217869 513770 217935 513773
rect 219390 513770 220064 513796
rect 217041 513768 220064 513770
rect 217041 513712 217046 513768
rect 217102 513712 217874 513768
rect 217930 513736 220064 513768
rect 396993 513770 397059 513773
rect 397126 513770 397132 513772
rect 396993 513768 397132 513770
rect 217930 513712 219450 513736
rect 217041 513710 219450 513712
rect 396993 513712 396998 513768
rect 397054 513712 397132 513768
rect 396993 513710 397132 513712
rect 217041 513707 217107 513710
rect 217869 513707 217935 513710
rect 396993 513707 397059 513710
rect 397126 513708 397132 513710
rect 397196 513770 397202 513772
rect 399342 513770 400016 513796
rect 397196 513736 400016 513770
rect 397196 513710 399402 513736
rect 397196 513708 397202 513710
rect 38009 513362 38075 513365
rect 38009 513360 40050 513362
rect 38009 513304 38014 513360
rect 38070 513304 40050 513360
rect 38009 513302 40050 513304
rect 38009 513299 38075 513302
rect 39990 512814 40050 513302
rect 217133 512818 217199 512821
rect 217685 512818 217751 512821
rect 219390 512818 220064 512844
rect 217133 512816 220064 512818
rect 217133 512760 217138 512816
rect 217194 512760 217690 512816
rect 217746 512784 220064 512816
rect 396625 512818 396691 512821
rect 396993 512818 397059 512821
rect 399342 512818 400016 512844
rect 396625 512816 400016 512818
rect 217746 512760 219450 512784
rect 217133 512758 219450 512760
rect 396625 512760 396630 512816
rect 396686 512760 396998 512816
rect 397054 512784 400016 512816
rect 397054 512760 399402 512784
rect 396625 512758 399402 512760
rect 217133 512755 217199 512758
rect 217685 512755 217751 512758
rect 396625 512755 396691 512758
rect 396993 512755 397059 512758
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 38101 511050 38167 511053
rect 217593 511050 217659 511053
rect 219390 511050 220064 511076
rect 38101 511048 40050 511050
rect 38101 510992 38106 511048
rect 38162 510992 40050 511048
rect 38101 510990 40050 510992
rect 217593 511048 220064 511050
rect 217593 510992 217598 511048
rect 217654 511016 220064 511048
rect 397085 511050 397151 511053
rect 399342 511050 400016 511076
rect 397085 511048 400016 511050
rect 217654 510992 219450 511016
rect 217593 510990 219450 510992
rect 397085 510992 397090 511048
rect 397146 511016 400016 511048
rect 397146 510992 399402 511016
rect 397085 510990 399402 510992
rect 38101 510987 38167 510990
rect 217593 510987 217659 510990
rect 397085 510987 397151 510990
rect 396901 510506 396967 510509
rect 397361 510506 397427 510509
rect 396901 510504 397427 510506
rect 396901 510448 396906 510504
rect 396962 510448 397366 510504
rect 397422 510448 397427 510504
rect 396901 510446 397427 510448
rect 396901 510443 396967 510446
rect 397361 510443 397427 510446
rect 38285 509962 38351 509965
rect 217501 509962 217567 509965
rect 219390 509962 220064 509988
rect 38285 509960 40050 509962
rect 38285 509904 38290 509960
rect 38346 509904 40050 509960
rect 38285 509902 40050 509904
rect 217501 509960 220064 509962
rect 217501 509904 217506 509960
rect 217562 509928 220064 509960
rect 396901 509962 396967 509965
rect 399342 509962 400016 509988
rect 396901 509960 400016 509962
rect 217562 509904 219450 509928
rect 217501 509902 219450 509904
rect 396901 509904 396906 509960
rect 396962 509928 400016 509960
rect 396962 509904 399402 509928
rect 396901 509902 399402 509904
rect 38285 509899 38351 509902
rect 217501 509899 217567 509902
rect 396901 509899 396967 509902
rect 217409 508194 217475 508197
rect 219390 508194 220064 508220
rect 217409 508192 220064 508194
rect 37825 507922 37891 507925
rect 38193 507922 38259 507925
rect 39990 507922 40050 508190
rect 217409 508136 217414 508192
rect 217470 508160 220064 508192
rect 396809 508194 396875 508197
rect 399342 508194 400016 508220
rect 396809 508192 400016 508194
rect 217470 508136 219450 508160
rect 217409 508134 219450 508136
rect 396809 508136 396814 508192
rect 396870 508160 400016 508192
rect 396870 508136 399402 508160
rect 396809 508134 399402 508136
rect 217409 508131 217475 508134
rect 396809 508131 396875 508134
rect 37825 507920 40050 507922
rect 37825 507864 37830 507920
rect 37886 507864 38198 507920
rect 38254 507864 40050 507920
rect 37825 507862 40050 507864
rect 37825 507859 37891 507862
rect 38193 507859 38259 507862
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 38561 489970 38627 489973
rect 217777 489970 217843 489973
rect 219390 489970 220064 489996
rect 38561 489968 40050 489970
rect 38561 489912 38566 489968
rect 38622 489912 40050 489968
rect 38561 489910 40050 489912
rect 217777 489968 220064 489970
rect 217777 489912 217782 489968
rect 217838 489936 220064 489968
rect 396717 489970 396783 489973
rect 399342 489970 400016 489996
rect 396717 489968 400016 489970
rect 217838 489912 219450 489936
rect 217777 489910 219450 489912
rect 396717 489912 396722 489968
rect 396778 489936 400016 489968
rect 396778 489912 399402 489936
rect 396717 489910 399402 489912
rect 38561 489907 38627 489910
rect 217777 489907 217843 489910
rect 396717 489907 396783 489910
rect -960 488596 480 488836
rect 37733 488338 37799 488341
rect 38326 488338 38332 488340
rect 37733 488336 38332 488338
rect 37733 488280 37738 488336
rect 37794 488280 38332 488336
rect 37733 488278 38332 488280
rect 37733 488275 37799 488278
rect 38326 488276 38332 488278
rect 38396 488338 38402 488340
rect 39438 488338 40020 488364
rect 38396 488304 40020 488338
rect 38396 488278 39498 488304
rect 38396 488276 38402 488278
rect 217910 488276 217916 488340
rect 217980 488338 217986 488340
rect 219390 488338 220064 488364
rect 217980 488304 220064 488338
rect 397177 488338 397243 488341
rect 399342 488338 400016 488364
rect 397177 488336 400016 488338
rect 217980 488278 219450 488304
rect 397177 488280 397182 488336
rect 397238 488304 400016 488336
rect 397238 488280 399402 488304
rect 397177 488278 399402 488280
rect 217980 488276 217986 488278
rect 397177 488275 397243 488278
rect 218421 488066 218487 488069
rect 219390 488066 220064 488092
rect 218421 488064 220064 488066
rect 38878 487460 38884 487524
rect 38948 487522 38954 487524
rect 39990 487522 40050 488062
rect 218421 488008 218426 488064
rect 218482 488032 220064 488064
rect 399342 488032 400016 488092
rect 218482 488008 219450 488032
rect 218421 488006 219450 488008
rect 218421 488003 218487 488006
rect 38948 487462 40050 487522
rect 38948 487460 38954 487462
rect 397177 487386 397243 487389
rect 397310 487386 397316 487388
rect 397177 487384 397316 487386
rect 397177 487328 397182 487384
rect 397238 487328 397316 487384
rect 397177 487326 397316 487328
rect 397177 487323 397243 487326
rect 397310 487324 397316 487326
rect 397380 487324 397386 487388
rect 180149 487250 180215 487253
rect 217910 487250 217916 487252
rect 180149 487248 217916 487250
rect 180149 487192 180154 487248
rect 180210 487192 217916 487248
rect 180149 487190 217916 487192
rect 180149 487187 180215 487190
rect 217910 487188 217916 487190
rect 217980 487188 217986 487252
rect 359406 487188 359412 487252
rect 359476 487250 359482 487252
rect 399342 487250 399402 488032
rect 359476 487190 399402 487250
rect 359476 487188 359482 487190
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 38469 480042 38535 480045
rect 217041 480042 217107 480045
rect 38469 480040 217107 480042
rect 38469 479984 38474 480040
rect 38530 479984 217046 480040
rect 217102 479984 217107 480040
rect 38469 479982 217107 479984
rect 38469 479979 38535 479982
rect 217041 479979 217107 479982
rect 56041 479636 56107 479637
rect 235993 479636 236059 479637
rect 56041 479632 56054 479636
rect 56118 479634 56124 479636
rect 235993 479634 236054 479636
rect 56041 479576 56046 479632
rect 56041 479572 56054 479576
rect 56118 479574 56198 479634
rect 235962 479632 236054 479634
rect 235962 479576 235998 479632
rect 235962 479574 236054 479576
rect 56118 479572 56124 479574
rect 235993 479572 236054 479574
rect 236118 479572 236124 479636
rect 56041 479571 56107 479572
rect 235993 479571 236059 479572
rect 217041 478954 217107 478957
rect 217174 478954 217180 478956
rect 217041 478952 217180 478954
rect 217041 478896 217046 478952
rect 217102 478896 217180 478952
rect 217041 478894 217180 478896
rect 217041 478891 217107 478894
rect 217174 478892 217180 478894
rect 217244 478892 217250 478956
rect 72325 478684 72391 478685
rect 74625 478684 74691 478685
rect 72325 478680 72372 478684
rect 72436 478682 72442 478684
rect 74574 478682 74580 478684
rect 72325 478624 72330 478680
rect 72325 478620 72372 478624
rect 72436 478622 72482 478682
rect 74534 478622 74580 478682
rect 74644 478680 74691 478684
rect 74686 478624 74691 478680
rect 72436 478620 72442 478622
rect 74574 478620 74580 478622
rect 74644 478620 74691 478624
rect 72325 478619 72391 478620
rect 74625 478619 74691 478620
rect 73153 478546 73219 478549
rect 76925 478548 76991 478549
rect 73470 478546 73476 478548
rect 73153 478544 73476 478546
rect 73153 478488 73158 478544
rect 73214 478488 73476 478544
rect 73153 478486 73476 478488
rect 73153 478483 73219 478486
rect 73470 478484 73476 478486
rect 73540 478484 73546 478548
rect 76925 478544 76972 478548
rect 77036 478546 77042 478548
rect 76925 478488 76930 478544
rect 76925 478484 76972 478488
rect 77036 478486 77082 478546
rect 77036 478484 77042 478486
rect 76925 478483 76991 478484
rect 75821 478412 75887 478413
rect 428549 478412 428615 478413
rect 430113 478412 430179 478413
rect 75821 478408 75868 478412
rect 75932 478410 75938 478412
rect 75821 478352 75826 478408
rect 75821 478348 75868 478352
rect 75932 478350 75978 478410
rect 428549 478408 428596 478412
rect 428660 478410 428666 478412
rect 430062 478410 430068 478412
rect 428549 478352 428554 478408
rect 75932 478348 75938 478350
rect 428549 478348 428596 478352
rect 428660 478350 428706 478410
rect 430022 478350 430068 478410
rect 430132 478408 430179 478412
rect 430174 478352 430179 478408
rect 428660 478348 428666 478350
rect 430062 478348 430068 478350
rect 430132 478348 430179 478352
rect 75821 478347 75887 478348
rect 428549 478347 428615 478348
rect 430113 478347 430179 478348
rect 79501 478276 79567 478277
rect 431309 478276 431375 478277
rect 432505 478276 432571 478277
rect 79501 478274 79548 478276
rect 79456 478272 79548 478274
rect 79456 478216 79506 478272
rect 79456 478214 79548 478216
rect 79501 478212 79548 478214
rect 79612 478212 79618 478276
rect 431309 478272 431356 478276
rect 431420 478274 431426 478276
rect 432454 478274 432460 478276
rect 431309 478216 431314 478272
rect 431309 478212 431356 478216
rect 431420 478214 431466 478274
rect 432414 478214 432460 478274
rect 432524 478272 432571 478276
rect 432566 478216 432571 478272
rect 431420 478212 431426 478214
rect 432454 478212 432460 478214
rect 432524 478212 432571 478216
rect 79501 478211 79567 478212
rect 431309 478211 431375 478212
rect 432505 478211 432571 478212
rect 80605 478140 80671 478141
rect 80605 478136 80652 478140
rect 80716 478138 80722 478140
rect 80605 478080 80610 478136
rect 80605 478076 80652 478080
rect 80716 478078 80762 478138
rect 80716 478076 80722 478078
rect 80605 478075 80671 478076
rect 86309 477596 86375 477597
rect 86309 477592 86356 477596
rect 86420 477594 86426 477596
rect 86309 477536 86314 477592
rect 86309 477532 86356 477536
rect 86420 477534 86466 477594
rect 86420 477532 86426 477534
rect 86309 477531 86375 477532
rect 63217 477460 63283 477461
rect 39798 477396 39804 477460
rect 39868 477458 39874 477460
rect 60590 477458 60596 477460
rect 39868 477398 60596 477458
rect 39868 477396 39874 477398
rect 60590 477396 60596 477398
rect 60660 477396 60666 477460
rect 63166 477458 63172 477460
rect 63126 477398 63172 477458
rect 63236 477456 63283 477460
rect 63278 477400 63283 477456
rect 63166 477396 63172 477398
rect 63236 477396 63283 477400
rect 63217 477395 63283 477396
rect 64229 477460 64295 477461
rect 64229 477456 64276 477460
rect 64340 477458 64346 477460
rect 64873 477458 64939 477461
rect 66529 477460 66595 477461
rect 67633 477460 67699 477461
rect 68737 477460 68803 477461
rect 70209 477460 70275 477461
rect 65374 477458 65380 477460
rect 64229 477400 64234 477456
rect 64229 477396 64276 477400
rect 64340 477398 64386 477458
rect 64873 477456 65380 477458
rect 64873 477400 64878 477456
rect 64934 477400 65380 477456
rect 64873 477398 65380 477400
rect 64340 477396 64346 477398
rect 64229 477395 64295 477396
rect 64873 477395 64939 477398
rect 65374 477396 65380 477398
rect 65444 477396 65450 477460
rect 66478 477458 66484 477460
rect 66438 477398 66484 477458
rect 66548 477456 66595 477460
rect 67582 477458 67588 477460
rect 66590 477400 66595 477456
rect 66478 477396 66484 477398
rect 66548 477396 66595 477400
rect 67542 477398 67588 477458
rect 67652 477456 67699 477460
rect 68686 477458 68692 477460
rect 67694 477400 67699 477456
rect 67582 477396 67588 477398
rect 67652 477396 67699 477400
rect 68646 477398 68692 477458
rect 68756 477456 68803 477460
rect 70158 477458 70164 477460
rect 68798 477400 68803 477456
rect 68686 477396 68692 477398
rect 68756 477396 68803 477400
rect 70118 477398 70164 477458
rect 70228 477456 70275 477460
rect 70270 477400 70275 477456
rect 70158 477396 70164 477398
rect 70228 477396 70275 477400
rect 66529 477395 66595 477396
rect 67633 477395 67699 477396
rect 68737 477395 68803 477396
rect 70209 477395 70275 477396
rect 70853 477458 70919 477461
rect 78121 477460 78187 477461
rect 71262 477458 71268 477460
rect 70853 477456 71268 477458
rect 70853 477400 70858 477456
rect 70914 477400 71268 477456
rect 70853 477398 71268 477400
rect 70853 477395 70919 477398
rect 71262 477396 71268 477398
rect 71332 477396 71338 477460
rect 78070 477458 78076 477460
rect 78030 477398 78076 477458
rect 78140 477456 78187 477460
rect 78182 477400 78187 477456
rect 78070 477396 78076 477398
rect 78140 477396 78187 477400
rect 81014 477396 81020 477460
rect 81084 477458 81090 477460
rect 81341 477458 81407 477461
rect 81801 477460 81867 477461
rect 81750 477458 81756 477460
rect 81084 477456 81407 477458
rect 81084 477400 81346 477456
rect 81402 477400 81407 477456
rect 81084 477398 81407 477400
rect 81710 477398 81756 477458
rect 81820 477456 81867 477460
rect 81862 477400 81867 477456
rect 81084 477396 81090 477398
rect 78121 477395 78187 477396
rect 81341 477395 81407 477398
rect 81750 477396 81756 477398
rect 81820 477396 81867 477400
rect 81801 477395 81867 477396
rect 82813 477460 82879 477461
rect 82813 477456 82860 477460
rect 82924 477458 82930 477460
rect 82813 477400 82818 477456
rect 82813 477396 82860 477400
rect 82924 477398 82970 477458
rect 82924 477396 82930 477398
rect 83590 477396 83596 477460
rect 83660 477458 83666 477460
rect 84101 477458 84167 477461
rect 85297 477460 85363 477461
rect 85246 477458 85252 477460
rect 83660 477456 84167 477458
rect 83660 477400 84106 477456
rect 84162 477400 84167 477456
rect 83660 477398 84167 477400
rect 85206 477398 85252 477458
rect 85316 477456 85363 477460
rect 85358 477400 85363 477456
rect 83660 477396 83666 477398
rect 82813 477395 82879 477396
rect 84101 477395 84167 477398
rect 85246 477396 85252 477398
rect 85316 477396 85363 477400
rect 85982 477396 85988 477460
rect 86052 477458 86058 477460
rect 86861 477458 86927 477461
rect 86052 477456 86927 477458
rect 86052 477400 86866 477456
rect 86922 477400 86927 477456
rect 86052 477398 86927 477400
rect 86052 477396 86058 477398
rect 85297 477395 85363 477396
rect 86861 477395 86927 477398
rect 87597 477460 87663 477461
rect 88241 477460 88307 477461
rect 87597 477456 87644 477460
rect 87708 477458 87714 477460
rect 87597 477400 87602 477456
rect 87597 477396 87644 477400
rect 87708 477398 87754 477458
rect 87708 477396 87714 477398
rect 88190 477396 88196 477460
rect 88260 477458 88307 477460
rect 88701 477460 88767 477461
rect 88260 477456 88352 477458
rect 88302 477400 88352 477456
rect 88260 477398 88352 477400
rect 88701 477456 88748 477460
rect 88812 477458 88818 477460
rect 89713 477458 89779 477461
rect 91185 477460 91251 477461
rect 89846 477458 89852 477460
rect 88701 477400 88706 477456
rect 88260 477396 88307 477398
rect 87597 477395 87663 477396
rect 88241 477395 88307 477396
rect 88701 477396 88748 477400
rect 88812 477398 88858 477458
rect 89713 477456 89852 477458
rect 89713 477400 89718 477456
rect 89774 477400 89852 477456
rect 89713 477398 89852 477400
rect 88812 477396 88818 477398
rect 88701 477395 88767 477396
rect 89713 477395 89779 477398
rect 89846 477396 89852 477398
rect 89916 477396 89922 477460
rect 91134 477458 91140 477460
rect 91094 477398 91140 477458
rect 91204 477456 91251 477460
rect 91246 477400 91251 477456
rect 91134 477396 91140 477398
rect 91204 477396 91251 477400
rect 91185 477395 91251 477396
rect 92197 477460 92263 477461
rect 92197 477456 92244 477460
rect 92308 477458 92314 477460
rect 93025 477458 93091 477461
rect 94405 477460 94471 477461
rect 95785 477460 95851 477461
rect 93342 477458 93348 477460
rect 92197 477400 92202 477456
rect 92197 477396 92244 477400
rect 92308 477398 92354 477458
rect 93025 477456 93348 477458
rect 93025 477400 93030 477456
rect 93086 477400 93348 477456
rect 93025 477398 93348 477400
rect 92308 477396 92314 477398
rect 92197 477395 92263 477396
rect 93025 477395 93091 477398
rect 93342 477396 93348 477398
rect 93412 477396 93418 477460
rect 94405 477456 94452 477460
rect 94516 477458 94522 477460
rect 95734 477458 95740 477460
rect 94405 477400 94410 477456
rect 94405 477396 94452 477400
rect 94516 477398 94562 477458
rect 95694 477398 95740 477458
rect 95804 477456 95851 477460
rect 95846 477400 95851 477456
rect 94516 477396 94522 477398
rect 95734 477396 95740 477398
rect 95804 477396 95851 477400
rect 94405 477395 94471 477396
rect 95785 477395 95851 477396
rect 96981 477460 97047 477461
rect 96981 477456 97028 477460
rect 97092 477458 97098 477460
rect 96981 477400 96986 477456
rect 96981 477396 97028 477400
rect 97092 477398 97138 477458
rect 97092 477396 97098 477398
rect 99046 477396 99052 477460
rect 99116 477458 99122 477460
rect 210693 477458 210759 477461
rect 219249 477458 219315 477461
rect 243169 477460 243235 477461
rect 244273 477460 244339 477461
rect 239622 477458 239628 477460
rect 99116 477456 210759 477458
rect 99116 477400 210698 477456
rect 210754 477400 210759 477456
rect 99116 477398 210759 477400
rect 99116 477396 99122 477398
rect 96981 477395 97047 477396
rect 210693 477395 210759 477398
rect 213134 477456 239628 477458
rect 213134 477400 219254 477456
rect 219310 477400 239628 477456
rect 213134 477398 239628 477400
rect 59445 477324 59511 477325
rect 59445 477320 59492 477324
rect 59556 477322 59562 477324
rect 60733 477322 60799 477325
rect 61694 477322 61700 477324
rect 59445 477264 59450 477320
rect 59445 477260 59492 477264
rect 59556 477262 59602 477322
rect 60733 477320 61700 477322
rect 60733 477264 60738 477320
rect 60794 477264 61700 477320
rect 60733 477262 61700 477264
rect 59556 477260 59562 477262
rect 59445 477259 59554 477260
rect 60733 477259 60799 477262
rect 61694 477260 61700 477262
rect 61764 477322 61770 477324
rect 210417 477322 210483 477325
rect 61764 477320 210483 477322
rect 61764 477264 210422 477320
rect 210478 477264 210483 477320
rect 61764 477262 210483 477264
rect 61764 477260 61770 477262
rect 210417 477259 210483 477262
rect 59494 477186 59554 477259
rect 210877 477186 210943 477189
rect 213134 477186 213194 477398
rect 219249 477395 219315 477398
rect 239622 477396 239628 477398
rect 239692 477396 239698 477460
rect 243118 477458 243124 477460
rect 243078 477398 243124 477458
rect 243188 477456 243235 477460
rect 244222 477458 244228 477460
rect 243230 477400 243235 477456
rect 243118 477396 243124 477398
rect 243188 477396 243235 477400
rect 244182 477398 244228 477458
rect 244292 477456 244339 477460
rect 244334 477400 244339 477456
rect 244222 477396 244228 477398
rect 244292 477396 244339 477400
rect 243169 477395 243235 477396
rect 244273 477395 244339 477396
rect 245469 477460 245535 477461
rect 245469 477456 245516 477460
rect 245580 477458 245586 477460
rect 245929 477458 245995 477461
rect 246430 477458 246436 477460
rect 245469 477400 245474 477456
rect 245469 477396 245516 477400
rect 245580 477398 245626 477458
rect 245929 477456 246436 477458
rect 245929 477400 245934 477456
rect 245990 477400 246436 477456
rect 245929 477398 246436 477400
rect 245580 477396 245586 477398
rect 245469 477395 245535 477396
rect 245929 477395 245995 477398
rect 246430 477396 246436 477398
rect 246500 477396 246506 477460
rect 247125 477458 247191 477461
rect 248597 477460 248663 477461
rect 250069 477460 250135 477461
rect 251265 477460 251331 477461
rect 252369 477460 252435 477461
rect 247534 477458 247540 477460
rect 247125 477456 247540 477458
rect 247125 477400 247130 477456
rect 247186 477400 247540 477456
rect 247125 477398 247540 477400
rect 247125 477395 247191 477398
rect 247534 477396 247540 477398
rect 247604 477396 247610 477460
rect 248597 477456 248644 477460
rect 248708 477458 248714 477460
rect 248597 477400 248602 477456
rect 248597 477396 248644 477400
rect 248708 477398 248754 477458
rect 250069 477456 250116 477460
rect 250180 477458 250186 477460
rect 251214 477458 251220 477460
rect 250069 477400 250074 477456
rect 248708 477396 248714 477398
rect 250069 477396 250116 477400
rect 250180 477398 250226 477458
rect 251174 477398 251220 477458
rect 251284 477456 251331 477460
rect 252318 477458 252324 477460
rect 251326 477400 251331 477456
rect 250180 477396 250186 477398
rect 251214 477396 251220 477398
rect 251284 477396 251331 477400
rect 252278 477398 252324 477458
rect 252388 477456 252435 477460
rect 252430 477400 252435 477456
rect 252318 477396 252324 477398
rect 252388 477396 252435 477400
rect 248597 477395 248663 477396
rect 250069 477395 250135 477396
rect 251265 477395 251331 477396
rect 252369 477395 252435 477396
rect 253381 477460 253447 477461
rect 254485 477460 254551 477461
rect 253381 477456 253428 477460
rect 253492 477458 253498 477460
rect 253381 477400 253386 477456
rect 253381 477396 253428 477400
rect 253492 477398 253538 477458
rect 254485 477456 254532 477460
rect 254596 477458 254602 477460
rect 255313 477458 255379 477461
rect 256969 477460 257035 477461
rect 260833 477460 260899 477461
rect 266353 477460 266419 477461
rect 255814 477458 255820 477460
rect 254485 477400 254490 477456
rect 253492 477396 253498 477398
rect 254485 477396 254532 477400
rect 254596 477398 254642 477458
rect 255313 477456 255820 477458
rect 255313 477400 255318 477456
rect 255374 477400 255820 477456
rect 255313 477398 255820 477400
rect 254596 477396 254602 477398
rect 253381 477395 253447 477396
rect 254485 477395 254551 477396
rect 255313 477395 255379 477398
rect 255814 477396 255820 477398
rect 255884 477396 255890 477460
rect 256918 477458 256924 477460
rect 256878 477398 256924 477458
rect 256988 477456 257035 477460
rect 260782 477458 260788 477460
rect 257030 477400 257035 477456
rect 256918 477396 256924 477398
rect 256988 477396 257035 477400
rect 260742 477398 260788 477458
rect 260852 477456 260899 477460
rect 260894 477400 260899 477456
rect 260782 477396 260788 477398
rect 260852 477396 260899 477400
rect 266302 477396 266308 477460
rect 266372 477458 266419 477460
rect 269113 477458 269179 477461
rect 269798 477458 269804 477460
rect 266372 477456 266464 477458
rect 266414 477400 266464 477456
rect 266372 477398 266464 477400
rect 269113 477456 269804 477458
rect 269113 477400 269118 477456
rect 269174 477400 269804 477456
rect 269113 477398 269804 477400
rect 266372 477396 266419 477398
rect 256969 477395 257035 477396
rect 260833 477395 260899 477396
rect 266353 477395 266419 477396
rect 269113 477395 269179 477398
rect 269798 477396 269804 477398
rect 269868 477396 269874 477460
rect 278773 477458 278839 477461
rect 279182 477458 279188 477460
rect 278773 477456 279188 477458
rect 278773 477400 278778 477456
rect 278834 477400 279188 477456
rect 278773 477398 279188 477400
rect 278773 477395 278839 477398
rect 279182 477396 279188 477398
rect 279252 477396 279258 477460
rect 415393 477458 415459 477461
rect 416078 477458 416084 477460
rect 415393 477456 416084 477458
rect 415393 477400 415398 477456
rect 415454 477400 416084 477456
rect 415393 477398 416084 477400
rect 415393 477395 415459 477398
rect 416078 477396 416084 477398
rect 416148 477396 416154 477460
rect 416773 477458 416839 477461
rect 417182 477458 417188 477460
rect 416773 477456 417188 477458
rect 416773 477400 416778 477456
rect 416834 477400 417188 477456
rect 416773 477398 417188 477400
rect 416773 477395 416839 477398
rect 417182 477396 417188 477398
rect 417252 477396 417258 477460
rect 418153 477458 418219 477461
rect 418286 477458 418292 477460
rect 418153 477456 418292 477458
rect 418153 477400 418158 477456
rect 418214 477400 418292 477456
rect 418153 477398 418292 477400
rect 418153 477395 418219 477398
rect 418286 477396 418292 477398
rect 418356 477396 418362 477460
rect 419533 477458 419599 477461
rect 420494 477458 420500 477460
rect 419533 477456 420500 477458
rect 419533 477400 419538 477456
rect 419594 477400 420500 477456
rect 419533 477398 420500 477400
rect 419533 477395 419599 477398
rect 420494 477396 420500 477398
rect 420564 477396 420570 477460
rect 420913 477458 420979 477461
rect 423121 477460 423187 477461
rect 421782 477458 421788 477460
rect 420913 477456 421788 477458
rect 420913 477400 420918 477456
rect 420974 477400 421788 477456
rect 420913 477398 421788 477400
rect 420913 477395 420979 477398
rect 421782 477396 421788 477398
rect 421852 477396 421858 477460
rect 423070 477458 423076 477460
rect 423030 477398 423076 477458
rect 423140 477456 423187 477460
rect 423182 477400 423187 477456
rect 423070 477396 423076 477398
rect 423140 477396 423187 477400
rect 423121 477395 423187 477396
rect 424133 477460 424199 477461
rect 425513 477460 425579 477461
rect 426617 477460 426683 477461
rect 427721 477460 427787 477461
rect 433425 477460 433491 477461
rect 434529 477460 434595 477461
rect 424133 477456 424180 477460
rect 424244 477458 424250 477460
rect 425462 477458 425468 477460
rect 424133 477400 424138 477456
rect 424133 477396 424180 477400
rect 424244 477398 424290 477458
rect 425422 477398 425468 477458
rect 425532 477456 425579 477460
rect 426566 477458 426572 477460
rect 425574 477400 425579 477456
rect 424244 477396 424250 477398
rect 425462 477396 425468 477398
rect 425532 477396 425579 477400
rect 426526 477398 426572 477458
rect 426636 477456 426683 477460
rect 427670 477458 427676 477460
rect 426678 477400 426683 477456
rect 426566 477396 426572 477398
rect 426636 477396 426683 477400
rect 427630 477398 427676 477458
rect 427740 477456 427787 477460
rect 433374 477458 433380 477460
rect 427782 477400 427787 477456
rect 427670 477396 427676 477398
rect 427740 477396 427787 477400
rect 433334 477398 433380 477458
rect 433444 477456 433491 477460
rect 434478 477458 434484 477460
rect 433486 477400 433491 477456
rect 433374 477396 433380 477398
rect 433444 477396 433491 477400
rect 434438 477398 434484 477458
rect 434548 477456 434595 477460
rect 434590 477400 434595 477456
rect 434478 477396 434484 477398
rect 434548 477396 434595 477400
rect 424133 477395 424199 477396
rect 425513 477395 425579 477396
rect 426617 477395 426683 477396
rect 427721 477395 427787 477396
rect 433425 477395 433491 477396
rect 434529 477395 434595 477396
rect 435725 477460 435791 477461
rect 435725 477456 435772 477460
rect 435836 477458 435842 477460
rect 436829 477458 436895 477461
rect 438117 477460 438183 477461
rect 437054 477458 437060 477460
rect 435725 477400 435730 477456
rect 435725 477396 435772 477400
rect 435836 477398 435882 477458
rect 436829 477456 437060 477458
rect 436829 477400 436834 477456
rect 436890 477400 437060 477456
rect 436829 477398 437060 477400
rect 435836 477396 435842 477398
rect 435725 477395 435791 477396
rect 436829 477395 436895 477398
rect 437054 477396 437060 477398
rect 437124 477396 437130 477460
rect 438117 477456 438164 477460
rect 438228 477458 438234 477460
rect 442993 477458 443059 477461
rect 443862 477458 443868 477460
rect 438117 477400 438122 477456
rect 438117 477396 438164 477400
rect 438228 477398 438274 477458
rect 442993 477456 443868 477458
rect 442993 477400 442998 477456
rect 443054 477400 443868 477456
rect 442993 477398 443868 477400
rect 438228 477396 438234 477398
rect 438117 477395 438183 477396
rect 442993 477395 443059 477398
rect 443862 477396 443868 477398
rect 443932 477396 443938 477460
rect 447133 477458 447199 477461
rect 447542 477458 447548 477460
rect 447133 477456 447548 477458
rect 447133 477400 447138 477456
rect 447194 477400 447548 477456
rect 447133 477398 447548 477400
rect 447133 477395 447199 477398
rect 447542 477396 447548 477398
rect 447612 477396 447618 477460
rect 448513 477458 448579 477461
rect 449750 477458 449756 477460
rect 448513 477456 449756 477458
rect 448513 477400 448518 477456
rect 448574 477400 449756 477456
rect 448513 477398 449756 477400
rect 448513 477395 448579 477398
rect 449750 477396 449756 477398
rect 449820 477396 449826 477460
rect 452653 477458 452719 477461
rect 453246 477458 453252 477460
rect 452653 477456 453252 477458
rect 452653 477400 452658 477456
rect 452714 477400 453252 477456
rect 452653 477398 453252 477400
rect 452653 477395 452719 477398
rect 453246 477396 453252 477398
rect 453316 477396 453322 477460
rect 213361 477322 213427 477325
rect 218881 477322 218947 477325
rect 237046 477322 237052 477324
rect 213361 477320 237052 477322
rect 213361 477264 213366 477320
rect 213422 477264 218886 477320
rect 218942 477264 237052 477320
rect 213361 477262 237052 477264
rect 213361 477259 213427 477262
rect 218881 477259 218947 477262
rect 237046 477260 237052 477262
rect 237116 477260 237122 477324
rect 258206 477260 258212 477324
rect 258276 477322 258282 477324
rect 259361 477322 259427 477325
rect 258276 477320 259427 477322
rect 258276 477264 259366 477320
rect 259422 477264 259427 477320
rect 258276 477262 259427 477264
rect 258276 477260 258282 477262
rect 259361 477259 259427 477262
rect 260833 477322 260899 477325
rect 261702 477322 261708 477324
rect 260833 477320 261708 477322
rect 260833 477264 260838 477320
rect 260894 477264 261708 477320
rect 260833 477262 261708 477264
rect 260833 477259 260899 477262
rect 261702 477260 261708 477262
rect 261772 477260 261778 477324
rect 263593 477322 263659 477325
rect 263910 477322 263916 477324
rect 263593 477320 263916 477322
rect 263593 477264 263598 477320
rect 263654 477264 263916 477320
rect 263593 477262 263916 477264
rect 263593 477259 263659 477262
rect 263910 477260 263916 477262
rect 263980 477260 263986 477324
rect 271873 477322 271939 477325
rect 272190 477322 272196 477324
rect 271873 477320 272196 477322
rect 271873 477264 271878 477320
rect 271934 477264 272196 477320
rect 271873 477262 272196 477264
rect 271873 477259 271939 477262
rect 272190 477260 272196 477262
rect 272260 477260 272266 477324
rect 276013 477322 276079 477325
rect 276974 477322 276980 477324
rect 276013 477320 276980 477322
rect 276013 477264 276018 477320
rect 276074 477264 276980 477320
rect 276013 477262 276980 477264
rect 276013 477259 276079 477262
rect 276974 477260 276980 477262
rect 277044 477260 277050 477324
rect 277669 477322 277735 477325
rect 278078 477322 278084 477324
rect 277669 477320 278084 477322
rect 277669 477264 277674 477320
rect 277730 477264 278084 477320
rect 277669 477262 278084 477264
rect 277669 477259 277735 477262
rect 278078 477260 278084 477262
rect 278148 477260 278154 477324
rect 398557 477322 398623 477325
rect 460974 477322 460980 477324
rect 398557 477320 460980 477322
rect 398557 477264 398562 477320
rect 398618 477264 460980 477320
rect 398557 477262 460980 477264
rect 398557 477259 398623 477262
rect 460974 477260 460980 477262
rect 461044 477260 461050 477324
rect 59494 477184 213194 477186
rect 59494 477128 210882 477184
rect 210938 477128 213194 477184
rect 59494 477126 213194 477128
rect 217501 477186 217567 477189
rect 217961 477186 218027 477189
rect 241646 477186 241652 477188
rect 217501 477184 241652 477186
rect 217501 477128 217506 477184
rect 217562 477128 217966 477184
rect 218022 477128 241652 477184
rect 217501 477126 241652 477128
rect 210877 477123 210943 477126
rect 217501 477123 217567 477126
rect 217961 477123 218027 477126
rect 241646 477124 241652 477126
rect 241716 477124 241722 477188
rect 273253 477186 273319 477189
rect 274398 477186 274404 477188
rect 273253 477184 274404 477186
rect 273253 477128 273258 477184
rect 273314 477128 274404 477184
rect 273253 477126 274404 477128
rect 273253 477123 273319 477126
rect 274398 477124 274404 477126
rect 274468 477124 274474 477188
rect 274633 477186 274699 477189
rect 275686 477186 275692 477188
rect 274633 477184 275692 477186
rect 274633 477128 274638 477184
rect 274694 477128 275692 477184
rect 274633 477126 275692 477128
rect 274633 477123 274699 477126
rect 275686 477124 275692 477126
rect 275756 477124 275762 477188
rect 311014 477124 311020 477188
rect 311084 477186 311090 477188
rect 311801 477186 311867 477189
rect 311084 477184 311867 477186
rect 311084 477128 311806 477184
rect 311862 477128 311867 477184
rect 311084 477126 311867 477128
rect 311084 477124 311090 477126
rect 311801 477123 311867 477126
rect 370497 477186 370563 477189
rect 435950 477186 435956 477188
rect 370497 477184 435956 477186
rect 370497 477128 370502 477184
rect 370558 477128 435956 477184
rect 370497 477126 435956 477128
rect 370497 477123 370563 477126
rect 435950 477124 435956 477126
rect 436020 477124 436026 477188
rect 438853 477186 438919 477189
rect 439446 477186 439452 477188
rect 438853 477184 439452 477186
rect 438853 477128 438858 477184
rect 438914 477128 439452 477184
rect 438853 477126 439452 477128
rect 438853 477123 438919 477126
rect 439446 477124 439452 477126
rect 439516 477186 439522 477188
rect 444189 477186 444255 477189
rect 439516 477184 444255 477186
rect 439516 477128 444194 477184
rect 444250 477128 444255 477184
rect 439516 477126 444255 477128
rect 439516 477124 439522 477126
rect 444189 477123 444255 477126
rect 444373 477186 444439 477189
rect 445334 477186 445340 477188
rect 444373 477184 445340 477186
rect 444373 477128 444378 477184
rect 444434 477128 445340 477184
rect 444373 477126 445340 477128
rect 444373 477123 444439 477126
rect 445334 477124 445340 477126
rect 445404 477124 445410 477188
rect 445753 477186 445819 477189
rect 446254 477186 446260 477188
rect 445753 477184 446260 477186
rect 445753 477128 445758 477184
rect 445814 477128 446260 477184
rect 445753 477126 446260 477128
rect 445753 477123 445819 477126
rect 446254 477124 446260 477126
rect 446324 477124 446330 477188
rect 448513 477186 448579 477189
rect 448646 477186 448652 477188
rect 448513 477184 448652 477186
rect 448513 477128 448518 477184
rect 448574 477128 448652 477184
rect 448513 477126 448652 477128
rect 448513 477123 448579 477126
rect 448646 477124 448652 477126
rect 448716 477124 448722 477188
rect 451365 477186 451431 477189
rect 452142 477186 452148 477188
rect 451365 477184 452148 477186
rect 451365 477128 451370 477184
rect 451426 477128 452148 477184
rect 451365 477126 452148 477128
rect 451365 477123 451431 477126
rect 452142 477124 452148 477126
rect 452212 477124 452218 477188
rect 458173 477186 458239 477189
rect 459134 477186 459140 477188
rect 458173 477184 459140 477186
rect 458173 477128 458178 477184
rect 458234 477128 459140 477184
rect 458173 477126 459140 477128
rect 458173 477123 458239 477126
rect 459134 477124 459140 477126
rect 459204 477124 459210 477188
rect 462313 477186 462379 477189
rect 463550 477186 463556 477188
rect 462313 477184 463556 477186
rect 462313 477128 462318 477184
rect 462374 477128 463556 477184
rect 462313 477126 463556 477128
rect 462313 477123 462379 477126
rect 463550 477124 463556 477126
rect 463620 477124 463626 477188
rect 60590 476988 60596 477052
rect 60660 477050 60666 477052
rect 213269 477050 213335 477053
rect 218973 477050 219039 477053
rect 240542 477050 240548 477052
rect 60660 477048 240548 477050
rect 60660 476992 213274 477048
rect 213330 476992 218978 477048
rect 219034 476992 240548 477048
rect 60660 476990 240548 476992
rect 60660 476988 60666 476990
rect 213269 476987 213335 476990
rect 218973 476987 219039 476990
rect 240542 476988 240548 476990
rect 240612 476988 240618 477052
rect 264973 477050 265039 477053
rect 265198 477050 265204 477052
rect 264973 477048 265204 477050
rect 264973 476992 264978 477048
rect 265034 476992 265204 477048
rect 264973 476990 265204 476992
rect 264973 476987 265039 476990
rect 265198 476988 265204 476990
rect 265268 476988 265274 477052
rect 270493 477050 270559 477053
rect 271270 477050 271276 477052
rect 270493 477048 271276 477050
rect 270493 476992 270498 477048
rect 270554 476992 271276 477048
rect 270493 476990 271276 476992
rect 270493 476987 270559 476990
rect 271270 476988 271276 476990
rect 271340 476988 271346 477052
rect 277577 477050 277643 477053
rect 278446 477050 278452 477052
rect 277577 477048 278452 477050
rect 277577 476992 277582 477048
rect 277638 476992 278452 477048
rect 277577 476990 278452 476992
rect 277577 476987 277643 476990
rect 278446 476988 278452 476990
rect 278516 476988 278522 477052
rect 285673 477050 285739 477053
rect 285990 477050 285996 477052
rect 285673 477048 285996 477050
rect 285673 476992 285678 477048
rect 285734 476992 285996 477048
rect 285673 476990 285996 476992
rect 285673 476987 285739 476990
rect 285990 476988 285996 476990
rect 286060 476988 286066 477052
rect 323342 476988 323348 477052
rect 323412 477050 323418 477052
rect 324221 477050 324287 477053
rect 323412 477048 324287 477050
rect 323412 476992 324226 477048
rect 324282 476992 324287 477048
rect 323412 476990 324287 476992
rect 323412 476988 323418 476990
rect 324221 476987 324287 476990
rect 325918 476988 325924 477052
rect 325988 477050 325994 477052
rect 326981 477050 327047 477053
rect 325988 477048 327047 477050
rect 325988 476992 326986 477048
rect 327042 476992 327047 477048
rect 325988 476990 327047 476992
rect 325988 476988 325994 476990
rect 326981 476987 327047 476990
rect 356881 477050 356947 477053
rect 438526 477050 438532 477052
rect 356881 477048 438532 477050
rect 356881 476992 356886 477048
rect 356942 476992 438532 477048
rect 356881 476990 438532 476992
rect 356881 476987 356947 476990
rect 438526 476988 438532 476990
rect 438596 476988 438602 477052
rect 440233 477050 440299 477053
rect 440734 477050 440740 477052
rect 440233 477048 440740 477050
rect 440233 476992 440238 477048
rect 440294 476992 440740 477048
rect 440233 476990 440740 476992
rect 440233 476987 440299 476990
rect 440734 476988 440740 476990
rect 440804 477050 440810 477052
rect 445661 477050 445727 477053
rect 440804 477048 445727 477050
rect 440804 476992 445666 477048
rect 445722 476992 445727 477048
rect 440804 476990 445727 476992
rect 440804 476988 440810 476990
rect 445661 476987 445727 476990
rect 446397 477050 446463 477053
rect 453614 477050 453620 477052
rect 446397 477048 453620 477050
rect 446397 476992 446402 477048
rect 446458 476992 453620 477048
rect 446397 476990 453620 476992
rect 446397 476987 446463 476990
rect 453614 476988 453620 476990
rect 453684 476988 453690 477052
rect 454033 477050 454099 477053
rect 454350 477050 454356 477052
rect 454033 477048 454356 477050
rect 454033 476992 454038 477048
rect 454094 476992 454356 477048
rect 454033 476990 454356 476992
rect 454033 476987 454099 476990
rect 454350 476988 454356 476990
rect 454420 476988 454426 477052
rect 456793 477050 456859 477053
rect 456926 477050 456932 477052
rect 456793 477048 456932 477050
rect 456793 476992 456798 477048
rect 456854 476992 456932 477048
rect 456793 476990 456932 476992
rect 456793 476987 456859 476990
rect 456926 476988 456932 476990
rect 456996 476988 457002 477052
rect 58157 476916 58223 476917
rect 58157 476914 58204 476916
rect 58076 476912 58204 476914
rect 58268 476914 58274 476916
rect 213177 476914 213243 476917
rect 219065 476914 219131 476917
rect 238150 476914 238156 476916
rect 58268 476912 238156 476914
rect 58076 476856 58162 476912
rect 58268 476856 213182 476912
rect 213238 476856 219070 476912
rect 219126 476856 238156 476912
rect 58076 476854 58204 476856
rect 58157 476852 58204 476854
rect 58268 476854 238156 476856
rect 58268 476852 58274 476854
rect 58157 476851 58223 476852
rect 213177 476851 213243 476854
rect 219065 476851 219131 476854
rect 238150 476852 238156 476854
rect 238220 476852 238226 476916
rect 255313 476914 255379 476917
rect 256182 476914 256188 476916
rect 255313 476912 256188 476914
rect 255313 476856 255318 476912
rect 255374 476856 256188 476912
rect 255313 476854 256188 476856
rect 255313 476851 255379 476854
rect 256182 476852 256188 476854
rect 256252 476852 256258 476916
rect 262213 476914 262279 476917
rect 262806 476914 262812 476916
rect 262213 476912 262812 476914
rect 262213 476856 262218 476912
rect 262274 476856 262812 476912
rect 262213 476854 262812 476856
rect 262213 476851 262279 476854
rect 262806 476852 262812 476854
rect 262876 476852 262882 476916
rect 270493 476914 270559 476917
rect 273253 476916 273319 476917
rect 270902 476914 270908 476916
rect 270493 476912 270908 476914
rect 270493 476856 270498 476912
rect 270554 476856 270908 476912
rect 270493 476854 270908 476856
rect 270493 476851 270559 476854
rect 270902 476852 270908 476854
rect 270972 476852 270978 476916
rect 273253 476914 273300 476916
rect 273208 476912 273300 476914
rect 273208 476856 273258 476912
rect 273208 476854 273300 476856
rect 273253 476852 273300 476854
rect 273364 476852 273370 476916
rect 320950 476852 320956 476916
rect 321020 476914 321026 476916
rect 321461 476914 321527 476917
rect 321020 476912 321527 476914
rect 321020 476856 321466 476912
rect 321522 476856 321527 476912
rect 321020 476854 321527 476856
rect 321020 476852 321026 476854
rect 273253 476851 273319 476852
rect 321461 476851 321527 476854
rect 357065 476914 357131 476917
rect 441613 476916 441679 476917
rect 441102 476914 441108 476916
rect 357065 476912 441108 476914
rect 357065 476856 357070 476912
rect 357126 476856 441108 476912
rect 357065 476854 441108 476856
rect 357065 476851 357131 476854
rect 441102 476852 441108 476854
rect 441172 476852 441178 476916
rect 441613 476912 441660 476916
rect 441724 476914 441730 476916
rect 455413 476914 455479 476917
rect 455638 476914 455644 476916
rect 441613 476856 441618 476912
rect 441613 476852 441660 476856
rect 441724 476854 441770 476914
rect 455413 476912 455644 476914
rect 455413 476856 455418 476912
rect 455474 476856 455644 476912
rect 455413 476854 455644 476856
rect 441724 476852 441730 476854
rect 441613 476851 441679 476852
rect 455413 476851 455479 476854
rect 455638 476852 455644 476854
rect 455708 476852 455714 476916
rect 456885 476914 456951 476917
rect 458030 476914 458036 476916
rect 456885 476912 458036 476914
rect 456885 476856 456890 476912
rect 456946 476856 458036 476912
rect 456885 476854 458036 476856
rect 456885 476851 456951 476854
rect 458030 476852 458036 476854
rect 458100 476852 458106 476916
rect 483013 476914 483079 476917
rect 483422 476914 483428 476916
rect 483013 476912 483428 476914
rect 483013 476856 483018 476912
rect 483074 476856 483428 476912
rect 483013 476854 483428 476856
rect 483013 476851 483079 476854
rect 483422 476852 483428 476854
rect 483492 476852 483498 476916
rect 57094 476716 57100 476780
rect 57164 476778 57170 476780
rect 57881 476778 57947 476781
rect 213361 476778 213427 476781
rect 57164 476776 213427 476778
rect 57164 476720 57886 476776
rect 57942 476720 213366 476776
rect 213422 476720 213427 476776
rect 57164 476718 213427 476720
rect 57164 476716 57170 476718
rect 57881 476715 57947 476718
rect 213361 476715 213427 476718
rect 266353 476778 266419 476781
rect 267590 476778 267596 476780
rect 266353 476776 267596 476778
rect 266353 476720 266358 476776
rect 266414 476720 267596 476776
rect 266353 476718 267596 476720
rect 266353 476715 266419 476718
rect 267590 476716 267596 476718
rect 267660 476716 267666 476780
rect 287697 476778 287763 476781
rect 288198 476778 288204 476780
rect 287697 476776 288204 476778
rect 287697 476720 287702 476776
rect 287758 476720 288204 476776
rect 287697 476718 288204 476720
rect 287697 476715 287763 476718
rect 288198 476716 288204 476718
rect 288268 476716 288274 476780
rect 300894 476716 300900 476780
rect 300964 476778 300970 476780
rect 302141 476778 302207 476781
rect 300964 476776 302207 476778
rect 300964 476720 302146 476776
rect 302202 476720 302207 476776
rect 300964 476718 302207 476720
rect 300964 476716 300970 476718
rect 302141 476715 302207 476718
rect 315798 476716 315804 476780
rect 315868 476778 315874 476780
rect 315941 476778 316007 476781
rect 315868 476776 316007 476778
rect 315868 476720 315946 476776
rect 316002 476720 316007 476776
rect 315868 476718 316007 476720
rect 315868 476716 315874 476718
rect 315941 476715 316007 476718
rect 318558 476716 318564 476780
rect 318628 476778 318634 476780
rect 318701 476778 318767 476781
rect 318628 476776 318767 476778
rect 318628 476720 318706 476776
rect 318762 476720 318767 476776
rect 318628 476718 318767 476720
rect 318628 476716 318634 476718
rect 318701 476715 318767 476718
rect 356697 476778 356763 476781
rect 456006 476778 456012 476780
rect 356697 476776 456012 476778
rect 356697 476720 356702 476776
rect 356758 476720 456012 476776
rect 356697 476718 456012 476720
rect 356697 476715 356763 476718
rect 456006 476716 456012 476718
rect 456076 476716 456082 476780
rect 490465 476778 490531 476781
rect 490966 476778 490972 476780
rect 490465 476776 490972 476778
rect 490465 476720 490470 476776
rect 490526 476720 490972 476776
rect 490465 476718 490972 476720
rect 490465 476715 490531 476718
rect 490966 476716 490972 476718
rect 491036 476716 491042 476780
rect 498193 476778 498259 476781
rect 498510 476778 498516 476780
rect 498193 476776 498516 476778
rect 498193 476720 498198 476776
rect 498254 476720 498516 476776
rect 498193 476718 498516 476720
rect 498193 476715 498259 476718
rect 498510 476716 498516 476718
rect 498580 476716 498586 476780
rect 84009 476644 84075 476645
rect 83958 476642 83964 476644
rect 83918 476582 83964 476642
rect 84028 476640 84075 476644
rect 210417 476642 210483 476645
rect 217501 476642 217567 476645
rect 259494 476642 259500 476644
rect 84070 476584 84075 476640
rect 83958 476580 83964 476582
rect 84028 476580 84075 476584
rect 84009 476579 84075 476580
rect 103470 476582 200130 476642
rect 91001 476508 91067 476509
rect 90950 476444 90956 476508
rect 91020 476506 91067 476508
rect 91020 476504 91112 476506
rect 91062 476448 91112 476504
rect 91020 476446 91112 476448
rect 91020 476444 91067 476446
rect 93526 476444 93532 476508
rect 93596 476506 93602 476508
rect 93761 476506 93827 476509
rect 93596 476504 93827 476506
rect 93596 476448 93766 476504
rect 93822 476448 93827 476504
rect 93596 476446 93827 476448
rect 93596 476444 93602 476446
rect 91001 476443 91067 476444
rect 93761 476443 93827 476446
rect 95969 476506 96035 476509
rect 99046 476506 99052 476508
rect 95969 476504 99052 476506
rect 95969 476448 95974 476504
rect 96030 476448 99052 476504
rect 95969 476446 99052 476448
rect 95969 476443 96035 476446
rect 99046 476444 99052 476446
rect 99116 476444 99122 476508
rect 79542 476308 79548 476372
rect 79612 476370 79618 476372
rect 98126 476370 98132 476372
rect 79612 476310 98132 476370
rect 79612 476308 79618 476310
rect 98126 476308 98132 476310
rect 98196 476370 98202 476372
rect 103470 476370 103530 476582
rect 200070 476506 200130 476582
rect 210417 476640 217567 476642
rect 210417 476584 210422 476640
rect 210478 476584 217506 476640
rect 217562 476584 217567 476640
rect 210417 476582 217567 476584
rect 210417 476579 210483 476582
rect 217501 476579 217567 476582
rect 217734 476582 259500 476642
rect 210509 476506 210575 476509
rect 214465 476506 214531 476509
rect 217734 476506 217794 476582
rect 259494 476580 259500 476582
rect 259564 476642 259570 476644
rect 263685 476642 263751 476645
rect 259564 476640 263751 476642
rect 259564 476584 263690 476640
rect 263746 476584 263751 476640
rect 259564 476582 263751 476584
rect 259564 476580 259570 476582
rect 263685 476579 263751 476582
rect 268193 476642 268259 476645
rect 268694 476642 268700 476644
rect 268193 476640 268700 476642
rect 268193 476584 268198 476640
rect 268254 476584 268700 476640
rect 268193 476582 268700 476584
rect 268193 476579 268259 476582
rect 268694 476580 268700 476582
rect 268764 476580 268770 476644
rect 308622 476580 308628 476644
rect 308692 476642 308698 476644
rect 309041 476642 309107 476645
rect 308692 476640 309107 476642
rect 308692 476584 309046 476640
rect 309102 476584 309107 476640
rect 308692 476582 309107 476584
rect 308692 476580 308698 476582
rect 309041 476579 309107 476582
rect 313406 476580 313412 476644
rect 313476 476642 313482 476644
rect 314561 476642 314627 476645
rect 313476 476640 314627 476642
rect 313476 476584 314566 476640
rect 314622 476584 314627 476640
rect 313476 476582 314627 476584
rect 313476 476580 313482 476582
rect 314561 476579 314627 476582
rect 398097 476642 398163 476645
rect 446397 476642 446463 476645
rect 398097 476640 446463 476642
rect 398097 476584 398102 476640
rect 398158 476584 446402 476640
rect 446458 476584 446463 476640
rect 398097 476582 446463 476584
rect 398097 476579 398163 476582
rect 446397 476579 446463 476582
rect 260782 476506 260788 476508
rect 200070 476504 217794 476506
rect 200070 476448 210514 476504
rect 210570 476448 214470 476504
rect 214526 476448 217794 476504
rect 200070 476446 217794 476448
rect 219390 476446 260788 476506
rect 210509 476443 210575 476446
rect 214465 476443 214531 476446
rect 98196 476310 103530 476370
rect 210693 476370 210759 476373
rect 214649 476370 214715 476373
rect 219390 476370 219450 476446
rect 260782 476444 260788 476446
rect 260852 476444 260858 476508
rect 289813 476506 289879 476509
rect 306097 476508 306163 476509
rect 290958 476506 290964 476508
rect 289813 476504 290964 476506
rect 289813 476448 289818 476504
rect 289874 476448 290964 476504
rect 289813 476446 290964 476448
rect 289813 476443 289879 476446
rect 290958 476444 290964 476446
rect 291028 476444 291034 476508
rect 306046 476444 306052 476508
rect 306116 476506 306163 476508
rect 419533 476508 419599 476509
rect 419533 476506 419580 476508
rect 306116 476504 306208 476506
rect 306158 476448 306208 476504
rect 306116 476446 306208 476448
rect 419488 476504 419580 476506
rect 419488 476448 419538 476504
rect 419488 476446 419580 476448
rect 306116 476444 306163 476446
rect 306097 476443 306163 476444
rect 419533 476444 419580 476446
rect 419644 476444 419650 476508
rect 433333 476506 433399 476509
rect 433742 476506 433748 476508
rect 433333 476504 433748 476506
rect 433333 476448 433338 476504
rect 433394 476448 433748 476504
rect 433333 476446 433748 476448
rect 419533 476443 419599 476444
rect 433333 476443 433399 476446
rect 433742 476444 433748 476446
rect 433812 476444 433818 476508
rect 441981 476506 442047 476509
rect 442758 476506 442764 476508
rect 441981 476504 442764 476506
rect 441981 476448 441986 476504
rect 442042 476448 442764 476504
rect 441981 476446 442764 476448
rect 441981 476443 442047 476446
rect 442758 476444 442764 476446
rect 442828 476444 442834 476508
rect 442993 476506 443059 476509
rect 443494 476506 443500 476508
rect 442993 476504 443500 476506
rect 442993 476448 442998 476504
rect 443054 476448 443500 476504
rect 442993 476446 443500 476448
rect 442993 476443 443059 476446
rect 443494 476444 443500 476446
rect 443564 476444 443570 476508
rect 449893 476506 449959 476509
rect 451038 476506 451044 476508
rect 449893 476504 451044 476506
rect 449893 476448 449898 476504
rect 449954 476448 451044 476504
rect 449893 476446 451044 476448
rect 449893 476443 449959 476446
rect 451038 476444 451044 476446
rect 451108 476444 451114 476508
rect 474733 476506 474799 476509
rect 475878 476506 475884 476508
rect 474733 476504 475884 476506
rect 474733 476448 474738 476504
rect 474794 476448 475884 476504
rect 474733 476446 475884 476448
rect 474733 476443 474799 476446
rect 475878 476444 475884 476446
rect 475948 476444 475954 476508
rect 477493 476506 477559 476509
rect 478454 476506 478460 476508
rect 477493 476504 478460 476506
rect 477493 476448 477498 476504
rect 477554 476448 478460 476504
rect 477493 476446 478460 476448
rect 477493 476443 477559 476446
rect 478454 476444 478460 476446
rect 478524 476444 478530 476508
rect 210693 476368 219450 476370
rect 210693 476312 210698 476368
rect 210754 476312 214654 476368
rect 214710 476312 219450 476368
rect 210693 476310 219450 476312
rect 98196 476308 98202 476310
rect 210693 476307 210759 476310
rect 214649 476307 214715 476310
rect 298502 476308 298508 476372
rect 298572 476370 298578 476372
rect 299381 476370 299447 476373
rect 303521 476372 303587 476373
rect 298572 476368 299447 476370
rect 298572 476312 299386 476368
rect 299442 476312 299447 476368
rect 298572 476310 299447 476312
rect 298572 476308 298578 476310
rect 299381 476307 299447 476310
rect 303470 476308 303476 476372
rect 303540 476370 303587 476372
rect 398281 476370 398347 476373
rect 458398 476370 458404 476372
rect 303540 476368 303632 476370
rect 303582 476312 303632 476368
rect 303540 476310 303632 476312
rect 398281 476368 458404 476370
rect 398281 476312 398286 476368
rect 398342 476312 458404 476368
rect 398281 476310 458404 476312
rect 303540 476308 303587 476310
rect 303521 476307 303587 476308
rect 398281 476307 398347 476310
rect 458398 476308 458404 476310
rect 458468 476308 458474 476372
rect 502333 476370 502399 476373
rect 503294 476370 503300 476372
rect 502333 476368 503300 476370
rect 502333 476312 502338 476368
rect 502394 476312 503300 476368
rect 502333 476310 503300 476312
rect 502333 476307 502399 476310
rect 503294 476308 503300 476310
rect 503364 476308 503370 476372
rect 68318 476172 68324 476236
rect 68388 476234 68394 476236
rect 68921 476234 68987 476237
rect 68388 476232 68987 476234
rect 68388 476176 68926 476232
rect 68982 476176 68987 476232
rect 68388 476174 68987 476176
rect 68388 476172 68394 476174
rect 68921 476171 68987 476174
rect 70710 476172 70716 476236
rect 70780 476234 70786 476236
rect 71681 476234 71747 476237
rect 70780 476232 71747 476234
rect 70780 476176 71686 476232
rect 71742 476176 71747 476232
rect 70780 476174 71747 476176
rect 70780 476172 70786 476174
rect 71681 476171 71747 476174
rect 73654 476172 73660 476236
rect 73724 476234 73730 476236
rect 74441 476234 74507 476237
rect 73724 476232 74507 476234
rect 73724 476176 74446 476232
rect 74502 476176 74507 476232
rect 73724 476174 74507 476176
rect 73724 476172 73730 476174
rect 74441 476171 74507 476174
rect 76046 476172 76052 476236
rect 76116 476234 76122 476236
rect 77201 476234 77267 476237
rect 76116 476232 77267 476234
rect 76116 476176 77206 476232
rect 77262 476176 77267 476232
rect 76116 476174 77267 476176
rect 76116 476172 76122 476174
rect 77201 476171 77267 476174
rect 78438 476172 78444 476236
rect 78508 476234 78514 476236
rect 78581 476234 78647 476237
rect 78508 476232 78647 476234
rect 78508 476176 78586 476232
rect 78642 476176 78647 476232
rect 78508 476174 78647 476176
rect 78508 476172 78514 476174
rect 78581 476171 78647 476174
rect 82721 476234 82787 476237
rect 95969 476234 96035 476237
rect 82721 476232 96035 476234
rect 82721 476176 82726 476232
rect 82782 476176 95974 476232
rect 96030 476176 96035 476232
rect 82721 476174 96035 476176
rect 82721 476171 82787 476174
rect 95969 476171 96035 476174
rect 96102 476172 96108 476236
rect 96172 476234 96178 476236
rect 96521 476234 96587 476237
rect 96172 476232 96587 476234
rect 96172 476176 96526 476232
rect 96582 476176 96587 476232
rect 96172 476174 96587 476176
rect 96172 476172 96178 476174
rect 96521 476171 96587 476174
rect 98494 476172 98500 476236
rect 98564 476234 98570 476236
rect 99281 476234 99347 476237
rect 98564 476232 99347 476234
rect 98564 476176 99286 476232
rect 99342 476176 99347 476232
rect 98564 476174 99347 476176
rect 98564 476172 98570 476174
rect 99281 476171 99347 476174
rect 100886 476172 100892 476236
rect 100956 476234 100962 476236
rect 102041 476234 102107 476237
rect 100956 476232 102107 476234
rect 100956 476176 102046 476232
rect 102102 476176 102107 476232
rect 100956 476174 102107 476176
rect 100956 476172 100962 476174
rect 102041 476171 102107 476174
rect 103646 476172 103652 476236
rect 103716 476234 103722 476236
rect 104801 476234 104867 476237
rect 103716 476232 104867 476234
rect 103716 476176 104806 476232
rect 104862 476176 104867 476232
rect 103716 476174 104867 476176
rect 103716 476172 103722 476174
rect 104801 476171 104867 476174
rect 106038 476172 106044 476236
rect 106108 476234 106114 476236
rect 106181 476234 106247 476237
rect 106108 476232 106247 476234
rect 106108 476176 106186 476232
rect 106242 476176 106247 476232
rect 106108 476174 106247 476176
rect 106108 476172 106114 476174
rect 106181 476171 106247 476174
rect 108246 476172 108252 476236
rect 108316 476234 108322 476236
rect 108941 476234 109007 476237
rect 108316 476232 109007 476234
rect 108316 476176 108946 476232
rect 109002 476176 109007 476232
rect 108316 476174 109007 476176
rect 108316 476172 108322 476174
rect 108941 476171 109007 476174
rect 111006 476172 111012 476236
rect 111076 476234 111082 476236
rect 111701 476234 111767 476237
rect 111076 476232 111767 476234
rect 111076 476176 111706 476232
rect 111762 476176 111767 476232
rect 111076 476174 111767 476176
rect 111076 476172 111082 476174
rect 111701 476171 111767 476174
rect 113398 476172 113404 476236
rect 113468 476234 113474 476236
rect 114461 476234 114527 476237
rect 113468 476232 114527 476234
rect 113468 476176 114466 476232
rect 114522 476176 114527 476232
rect 113468 476174 114527 476176
rect 113468 476172 113474 476174
rect 114461 476171 114527 476174
rect 115974 476172 115980 476236
rect 116044 476234 116050 476236
rect 117221 476234 117287 476237
rect 118601 476236 118667 476237
rect 116044 476232 117287 476234
rect 116044 476176 117226 476232
rect 117282 476176 117287 476232
rect 116044 476174 117287 476176
rect 116044 476172 116050 476174
rect 117221 476171 117287 476174
rect 118550 476172 118556 476236
rect 118620 476234 118667 476236
rect 118620 476232 118712 476234
rect 118662 476176 118712 476232
rect 118620 476174 118712 476176
rect 118620 476172 118667 476174
rect 120942 476172 120948 476236
rect 121012 476234 121018 476236
rect 121361 476234 121427 476237
rect 121012 476232 121427 476234
rect 121012 476176 121366 476232
rect 121422 476176 121427 476232
rect 121012 476174 121427 476176
rect 121012 476172 121018 476174
rect 118601 476171 118667 476172
rect 121361 476171 121427 476174
rect 123518 476172 123524 476236
rect 123588 476234 123594 476236
rect 124121 476234 124187 476237
rect 123588 476232 124187 476234
rect 123588 476176 124126 476232
rect 124182 476176 124187 476232
rect 123588 476174 124187 476176
rect 123588 476172 123594 476174
rect 124121 476171 124187 476174
rect 125910 476172 125916 476236
rect 125980 476234 125986 476236
rect 126881 476234 126947 476237
rect 125980 476232 126947 476234
rect 125980 476176 126886 476232
rect 126942 476176 126947 476232
rect 125980 476174 126947 476176
rect 125980 476172 125986 476174
rect 126881 476171 126947 476174
rect 128486 476172 128492 476236
rect 128556 476234 128562 476236
rect 129641 476234 129707 476237
rect 131021 476236 131087 476237
rect 131021 476234 131068 476236
rect 128556 476232 129707 476234
rect 128556 476176 129646 476232
rect 129702 476176 129707 476232
rect 128556 476174 129707 476176
rect 130976 476232 131068 476234
rect 130976 476176 131026 476232
rect 130976 476174 131068 476176
rect 128556 476172 128562 476174
rect 129641 476171 129707 476174
rect 131021 476172 131068 476174
rect 131132 476172 131138 476236
rect 133454 476172 133460 476236
rect 133524 476234 133530 476236
rect 133781 476234 133847 476237
rect 133524 476232 133847 476234
rect 133524 476176 133786 476232
rect 133842 476176 133847 476232
rect 133524 476174 133847 476176
rect 133524 476172 133530 476174
rect 131021 476171 131087 476172
rect 133781 476171 133847 476174
rect 135846 476172 135852 476236
rect 135916 476234 135922 476236
rect 136541 476234 136607 476237
rect 135916 476232 136607 476234
rect 135916 476176 136546 476232
rect 136602 476176 136607 476232
rect 135916 476174 136607 476176
rect 135916 476172 135922 476174
rect 136541 476171 136607 476174
rect 138422 476172 138428 476236
rect 138492 476234 138498 476236
rect 139301 476234 139367 476237
rect 138492 476232 139367 476234
rect 138492 476176 139306 476232
rect 139362 476176 139367 476232
rect 138492 476174 139367 476176
rect 138492 476172 138498 476174
rect 139301 476171 139367 476174
rect 140998 476172 141004 476236
rect 141068 476234 141074 476236
rect 142061 476234 142127 476237
rect 143441 476236 143507 476237
rect 141068 476232 142127 476234
rect 141068 476176 142066 476232
rect 142122 476176 142127 476232
rect 141068 476174 142127 476176
rect 141068 476172 141074 476174
rect 142061 476171 142127 476174
rect 143390 476172 143396 476236
rect 143460 476234 143507 476236
rect 143460 476232 143552 476234
rect 143502 476176 143552 476232
rect 143460 476174 143552 476176
rect 143460 476172 143507 476174
rect 145966 476172 145972 476236
rect 146036 476234 146042 476236
rect 146201 476234 146267 476237
rect 146036 476232 146267 476234
rect 146036 476176 146206 476232
rect 146262 476176 146267 476232
rect 146036 476174 146267 476176
rect 146036 476172 146042 476174
rect 143441 476171 143507 476172
rect 146201 476171 146267 476174
rect 247033 476234 247099 476237
rect 248270 476234 248276 476236
rect 247033 476232 248276 476234
rect 247033 476176 247038 476232
rect 247094 476176 248276 476232
rect 247033 476174 248276 476176
rect 247033 476171 247099 476174
rect 248270 476172 248276 476174
rect 248340 476172 248346 476236
rect 249793 476234 249859 476237
rect 250662 476234 250668 476236
rect 249793 476232 250668 476234
rect 249793 476176 249798 476232
rect 249854 476176 250668 476232
rect 249793 476174 250668 476176
rect 249793 476171 249859 476174
rect 250662 476172 250668 476174
rect 250732 476172 250738 476236
rect 252553 476234 252619 476237
rect 253606 476234 253612 476236
rect 252553 476232 253612 476234
rect 252553 476176 252558 476232
rect 252614 476176 253612 476232
rect 252553 476174 253612 476176
rect 252553 476171 252619 476174
rect 253606 476172 253612 476174
rect 253676 476172 253682 476236
rect 258257 476234 258323 476237
rect 258390 476234 258396 476236
rect 258257 476232 258396 476234
rect 258257 476176 258262 476232
rect 258318 476176 258396 476232
rect 258257 476174 258396 476176
rect 258257 476171 258323 476174
rect 258390 476172 258396 476174
rect 258460 476172 258466 476236
rect 260833 476234 260899 476237
rect 263593 476236 263659 476237
rect 260966 476234 260972 476236
rect 260833 476232 260972 476234
rect 260833 476176 260838 476232
rect 260894 476176 260972 476232
rect 260833 476174 260972 476176
rect 260833 476171 260899 476174
rect 260966 476172 260972 476174
rect 261036 476172 261042 476236
rect 263542 476172 263548 476236
rect 263612 476234 263659 476236
rect 264973 476234 265039 476237
rect 265934 476234 265940 476236
rect 263612 476232 263704 476234
rect 263654 476176 263704 476232
rect 263612 476174 263704 476176
rect 264973 476232 265940 476234
rect 264973 476176 264978 476232
rect 265034 476176 265940 476232
rect 264973 476174 265940 476176
rect 263612 476172 263659 476174
rect 263593 476171 263659 476172
rect 264973 476171 265039 476174
rect 265934 476172 265940 476174
rect 266004 476172 266010 476236
rect 268009 476234 268075 476237
rect 268326 476234 268332 476236
rect 268009 476232 268332 476234
rect 268009 476176 268014 476232
rect 268070 476176 268332 476232
rect 268009 476174 268332 476176
rect 268009 476171 268075 476174
rect 268326 476172 268332 476174
rect 268396 476172 268402 476236
rect 273253 476234 273319 476237
rect 276013 476236 276079 476237
rect 273478 476234 273484 476236
rect 273253 476232 273484 476234
rect 273253 476176 273258 476232
rect 273314 476176 273484 476232
rect 273253 476174 273484 476176
rect 273253 476171 273319 476174
rect 273478 476172 273484 476174
rect 273548 476172 273554 476236
rect 276013 476234 276060 476236
rect 275968 476232 276060 476234
rect 275968 476176 276018 476232
rect 275968 476174 276060 476176
rect 276013 476172 276060 476174
rect 276124 476172 276130 476236
rect 280153 476234 280219 476237
rect 280838 476234 280844 476236
rect 280153 476232 280844 476234
rect 280153 476176 280158 476232
rect 280214 476176 280844 476232
rect 280153 476174 280844 476176
rect 276013 476171 276079 476172
rect 280153 476171 280219 476174
rect 280838 476172 280844 476174
rect 280908 476172 280914 476236
rect 282913 476234 282979 476237
rect 283414 476234 283420 476236
rect 282913 476232 283420 476234
rect 282913 476176 282918 476232
rect 282974 476176 283420 476232
rect 282913 476174 283420 476176
rect 282913 476171 282979 476174
rect 283414 476172 283420 476174
rect 283484 476172 283490 476236
rect 292573 476234 292639 476237
rect 293350 476234 293356 476236
rect 292573 476232 293356 476234
rect 292573 476176 292578 476232
rect 292634 476176 293356 476232
rect 292573 476174 293356 476176
rect 292573 476171 292639 476174
rect 293350 476172 293356 476174
rect 293420 476172 293426 476236
rect 295926 476172 295932 476236
rect 295996 476234 296002 476236
rect 296253 476234 296319 476237
rect 295996 476232 296319 476234
rect 295996 476176 296258 476232
rect 296314 476176 296319 476232
rect 295996 476174 296319 476176
rect 295996 476172 296002 476174
rect 296253 476171 296319 476174
rect 427813 476234 427879 476237
rect 430573 476236 430639 476237
rect 428222 476234 428228 476236
rect 427813 476232 428228 476234
rect 427813 476176 427818 476232
rect 427874 476176 428228 476232
rect 427813 476174 428228 476176
rect 427813 476171 427879 476174
rect 428222 476172 428228 476174
rect 428292 476172 428298 476236
rect 430573 476234 430620 476236
rect 430528 476232 430620 476234
rect 430528 476176 430578 476232
rect 430528 476174 430620 476176
rect 430573 476172 430620 476174
rect 430684 476172 430690 476236
rect 445753 476234 445819 476237
rect 445886 476234 445892 476236
rect 445753 476232 445892 476234
rect 445753 476176 445758 476232
rect 445814 476176 445892 476232
rect 445753 476174 445892 476176
rect 430573 476171 430639 476172
rect 445753 476171 445819 476174
rect 445886 476172 445892 476174
rect 445956 476172 445962 476236
rect 447133 476234 447199 476237
rect 448278 476234 448284 476236
rect 447133 476232 448284 476234
rect 447133 476176 447138 476232
rect 447194 476176 448284 476232
rect 447133 476174 448284 476176
rect 447133 476171 447199 476174
rect 448278 476172 448284 476174
rect 448348 476172 448354 476236
rect 449893 476234 449959 476237
rect 450854 476234 450860 476236
rect 449893 476232 450860 476234
rect 449893 476176 449898 476232
rect 449954 476176 450860 476232
rect 449893 476174 450860 476176
rect 449893 476171 449959 476174
rect 450854 476172 450860 476174
rect 450924 476172 450930 476236
rect 465073 476234 465139 476237
rect 465942 476234 465948 476236
rect 465073 476232 465948 476234
rect 465073 476176 465078 476232
rect 465134 476176 465948 476232
rect 465073 476174 465948 476176
rect 465073 476171 465139 476174
rect 465942 476172 465948 476174
rect 466012 476172 466018 476236
rect 467833 476234 467899 476237
rect 468150 476234 468156 476236
rect 467833 476232 468156 476234
rect 467833 476176 467838 476232
rect 467894 476176 468156 476232
rect 467833 476174 468156 476176
rect 467833 476171 467899 476174
rect 468150 476172 468156 476174
rect 468220 476172 468226 476236
rect 470777 476234 470843 476237
rect 470910 476234 470916 476236
rect 470777 476232 470916 476234
rect 470777 476176 470782 476232
rect 470838 476176 470916 476232
rect 470777 476174 470916 476176
rect 470777 476171 470843 476174
rect 470910 476172 470916 476174
rect 470980 476172 470986 476236
rect 473353 476234 473419 476237
rect 473486 476234 473492 476236
rect 473353 476232 473492 476234
rect 473353 476176 473358 476232
rect 473414 476176 473492 476232
rect 473353 476174 473492 476176
rect 473353 476171 473419 476174
rect 473486 476172 473492 476174
rect 473556 476172 473562 476236
rect 480529 476234 480595 476237
rect 480846 476234 480852 476236
rect 480529 476232 480852 476234
rect 480529 476176 480534 476232
rect 480590 476176 480852 476232
rect 480529 476174 480852 476176
rect 480529 476171 480595 476174
rect 480846 476172 480852 476174
rect 480916 476172 480922 476236
rect 485773 476234 485839 476237
rect 488533 476236 488599 476237
rect 485998 476234 486004 476236
rect 485773 476232 486004 476234
rect 485773 476176 485778 476232
rect 485834 476176 486004 476232
rect 485773 476174 486004 476176
rect 485773 476171 485839 476174
rect 485998 476172 486004 476174
rect 486068 476172 486074 476236
rect 488533 476234 488580 476236
rect 488488 476232 488580 476234
rect 488488 476176 488538 476232
rect 488488 476174 488580 476176
rect 488533 476172 488580 476174
rect 488644 476172 488650 476236
rect 492673 476234 492739 476237
rect 493358 476234 493364 476236
rect 492673 476232 493364 476234
rect 492673 476176 492678 476232
rect 492734 476176 493364 476232
rect 492673 476174 493364 476176
rect 488533 476171 488599 476172
rect 492673 476171 492739 476174
rect 493358 476172 493364 476174
rect 493428 476172 493434 476236
rect 495433 476234 495499 476237
rect 500953 476236 501019 476237
rect 495934 476234 495940 476236
rect 495433 476232 495940 476234
rect 495433 476176 495438 476232
rect 495494 476176 495940 476232
rect 495433 476174 495940 476176
rect 495433 476171 495499 476174
rect 495934 476172 495940 476174
rect 496004 476172 496010 476236
rect 500902 476172 500908 476236
rect 500972 476234 501019 476236
rect 505093 476234 505159 476237
rect 505870 476234 505876 476236
rect 500972 476232 501064 476234
rect 501014 476176 501064 476232
rect 500972 476174 501064 476176
rect 505093 476232 505876 476234
rect 505093 476176 505098 476232
rect 505154 476176 505876 476232
rect 505093 476174 505876 476176
rect 500972 476172 501019 476174
rect 500953 476171 501019 476172
rect 505093 476171 505159 476174
rect 505870 476172 505876 476174
rect 505940 476172 505946 476236
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 217726 474676 217732 474740
rect 217796 474738 217802 474740
rect 218145 474738 218211 474741
rect 217796 474736 218211 474738
rect 217796 474680 218150 474736
rect 218206 474680 218211 474736
rect 217796 474678 218211 474680
rect 217796 474676 217802 474678
rect 218145 474675 218211 474678
rect 218830 474676 218836 474740
rect 218900 474738 218906 474740
rect 219893 474738 219959 474741
rect 218900 474736 219959 474738
rect 218900 474680 219898 474736
rect 219954 474680 219959 474736
rect 218900 474678 219959 474680
rect 218900 474676 218906 474678
rect 219893 474675 219959 474678
rect 399518 474540 399524 474604
rect 399588 474602 399594 474604
rect 442993 474602 443059 474605
rect 399588 474600 443059 474602
rect 399588 474544 442998 474600
rect 443054 474544 443059 474600
rect 399588 474542 443059 474544
rect 399588 474540 399594 474542
rect 442993 474539 443059 474542
rect 398189 474466 398255 474469
rect 462313 474466 462379 474469
rect 398189 474464 462379 474466
rect 398189 474408 398194 474464
rect 398250 474408 462318 474464
rect 462374 474408 462379 474464
rect 398189 474406 462379 474408
rect 398189 474403 398255 474406
rect 462313 474403 462379 474406
rect 397821 474330 397887 474333
rect 467833 474330 467899 474333
rect 397821 474328 467899 474330
rect 397821 474272 397826 474328
rect 397882 474272 467838 474328
rect 467894 474272 467899 474328
rect 397821 474270 467899 474272
rect 397821 474267 397887 474270
rect 467833 474267 467899 474270
rect 218881 474194 218947 474197
rect 255313 474194 255379 474197
rect 218881 474192 255379 474194
rect 218881 474136 218886 474192
rect 218942 474136 255318 474192
rect 255374 474136 255379 474192
rect 218881 474134 255379 474136
rect 218881 474131 218947 474134
rect 255313 474131 255379 474134
rect 398465 474194 398531 474197
rect 470777 474194 470843 474197
rect 398465 474192 470843 474194
rect 398465 474136 398470 474192
rect 398526 474136 470782 474192
rect 470838 474136 470843 474192
rect 398465 474134 470843 474136
rect 398465 474131 398531 474134
rect 470777 474131 470843 474134
rect 216121 474058 216187 474061
rect 258257 474058 258323 474061
rect 216121 474056 258323 474058
rect 216121 474000 216126 474056
rect 216182 474000 258262 474056
rect 258318 474000 258323 474056
rect 216121 473998 258323 474000
rect 216121 473995 216187 473998
rect 258257 473995 258323 473998
rect 398005 474058 398071 474061
rect 473353 474058 473419 474061
rect 398005 474056 473419 474058
rect 398005 474000 398010 474056
rect 398066 474000 473358 474056
rect 473414 474000 473419 474056
rect 398005 473998 473419 474000
rect 398005 473995 398071 473998
rect 473353 473995 473419 473998
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 216070 461484 216076 461548
rect 216140 461546 216146 461548
rect 430573 461546 430639 461549
rect 216140 461544 430639 461546
rect 216140 461488 430578 461544
rect 430634 461488 430639 461544
rect 216140 461486 430639 461488
rect 216140 461484 216146 461486
rect 430573 461483 430639 461486
rect 212206 460124 212212 460188
rect 212276 460186 212282 460188
rect 427813 460186 427879 460189
rect 212276 460184 427879 460186
rect 212276 460128 427818 460184
rect 427874 460128 427879 460184
rect 212276 460126 427879 460128
rect 212276 460124 212282 460126
rect 427813 460123 427879 460126
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 397310 446388 397316 446452
rect 397380 446450 397386 446452
rect 530485 446450 530551 446453
rect 530894 446450 530900 446452
rect 397380 446448 530900 446450
rect 397380 446392 530490 446448
rect 530546 446392 530900 446448
rect 397380 446390 530900 446392
rect 397380 446388 397386 446390
rect 530485 446387 530551 446390
rect 530894 446388 530900 446390
rect 530964 446388 530970 446452
rect 170857 445772 170923 445773
rect 170806 445770 170812 445772
rect 170766 445710 170812 445770
rect 170876 445768 170923 445772
rect 170918 445712 170923 445768
rect 170806 445708 170812 445710
rect 170876 445708 170923 445712
rect 350942 445708 350948 445772
rect 351012 445770 351018 445772
rect 351085 445770 351151 445773
rect 351012 445768 351151 445770
rect 351012 445712 351090 445768
rect 351146 445712 351151 445768
rect 351012 445710 351151 445712
rect 351012 445708 351018 445710
rect 170857 445707 170923 445708
rect 351085 445707 351151 445710
rect 111701 445226 111767 445229
rect 214782 445226 214788 445228
rect 111701 445224 214788 445226
rect 111701 445168 111706 445224
rect 111762 445168 214788 445224
rect 111701 445166 214788 445168
rect 111701 445163 111767 445166
rect 214782 445164 214788 445166
rect 214852 445164 214858 445228
rect 108941 445090 109007 445093
rect 214598 445090 214604 445092
rect 108941 445088 214604 445090
rect 108941 445032 108946 445088
rect 109002 445032 214604 445088
rect 108941 445030 214604 445032
rect 108941 445027 109007 445030
rect 214598 445028 214604 445030
rect 214668 445028 214674 445092
rect 93761 444954 93827 444957
rect 216806 444954 216812 444956
rect 93761 444952 216812 444954
rect 93761 444896 93766 444952
rect 93822 444896 216812 444952
rect 93761 444894 216812 444896
rect 93761 444891 93827 444894
rect 216806 444892 216812 444894
rect 216876 444892 216882 444956
rect 583520 444668 584960 444908
rect 398782 444212 398788 444276
rect 398852 444274 398858 444276
rect 400121 444274 400187 444277
rect 398852 444272 400187 444274
rect 398852 444216 400126 444272
rect 400182 444216 400187 444272
rect 398852 444214 400187 444216
rect 398852 444212 398858 444214
rect 400121 444211 400187 444214
rect 74441 443594 74507 443597
rect 216622 443594 216628 443596
rect 74441 443592 216628 443594
rect 74441 443536 74446 443592
rect 74502 443536 216628 443592
rect 74441 443534 216628 443536
rect 74441 443531 74507 443534
rect 216622 443532 216628 443534
rect 216692 443532 216698 443596
rect 538213 439786 538279 439789
rect 536558 439784 538279 439786
rect 536558 439728 538218 439784
rect 538274 439728 538279 439784
rect 536558 439726 538279 439728
rect 178493 439242 178559 439245
rect 358813 439242 358879 439245
rect 177070 439240 178559 439242
rect 177070 439220 178498 439240
rect 176548 439184 178498 439220
rect 178554 439184 178559 439240
rect 176548 439182 178559 439184
rect 356562 439240 358879 439242
rect 356562 439184 358818 439240
rect 358874 439184 358879 439240
rect 536558 439190 536618 439726
rect 538213 439723 538279 439726
rect 356562 439182 358879 439184
rect 176548 439160 177130 439182
rect 178493 439179 178559 439182
rect 358813 439179 358879 439182
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580441 418298 580507 418301
rect 583520 418298 584960 418388
rect 580441 418296 584960 418298
rect 580441 418240 580446 418296
rect 580502 418240 584960 418296
rect 580441 418238 584960 418240
rect 580441 418235 580507 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3509 410546 3575 410549
rect -960 410544 3575 410546
rect -960 410488 3514 410544
rect 3570 410488 3575 410544
rect -960 410486 3575 410488
rect -960 410396 480 410486
rect 3509 410483 3575 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 38469 397354 38535 397357
rect 38469 397352 40050 397354
rect 38469 397296 38474 397352
rect 38530 397296 40050 397352
rect 38469 397294 40050 397296
rect 38469 397291 38535 397294
rect 39990 396894 40050 397294
rect 217685 396946 217751 396949
rect 396625 396946 396691 396949
rect 217685 396944 219450 396946
rect 217685 396888 217690 396944
rect 217746 396924 219450 396944
rect 396625 396944 399402 396946
rect 217746 396888 220064 396924
rect 217685 396886 220064 396888
rect 217685 396883 217751 396886
rect 219390 396864 220064 396886
rect 396625 396888 396630 396944
rect 396686 396924 399402 396944
rect 396686 396888 400016 396924
rect 396625 396886 400016 396888
rect 396625 396883 396691 396886
rect 399342 396864 400016 396886
rect 217317 395994 217383 395997
rect 218789 395994 218855 395997
rect 396533 395994 396599 395997
rect 217317 395992 219450 395994
rect 38469 395450 38535 395453
rect 39990 395450 40050 395942
rect 217317 395936 217322 395992
rect 217378 395936 218794 395992
rect 218850 395972 219450 395992
rect 396533 395992 399402 395994
rect 218850 395936 220064 395972
rect 217317 395934 220064 395936
rect 217317 395931 217383 395934
rect 218789 395931 218855 395934
rect 219390 395912 220064 395934
rect 396533 395936 396538 395992
rect 396594 395972 399402 395992
rect 396594 395936 400016 395972
rect 396533 395934 400016 395936
rect 396533 395931 396599 395934
rect 399342 395912 400016 395934
rect 38469 395448 40050 395450
rect 38469 395392 38474 395448
rect 38530 395392 40050 395448
rect 38469 395390 40050 395392
rect 38469 395387 38535 395390
rect 396625 394634 396691 394637
rect 397126 394634 397132 394636
rect 396625 394632 397132 394634
rect 396625 394576 396630 394632
rect 396686 394576 397132 394632
rect 396625 394574 397132 394576
rect 396625 394571 396691 394574
rect 397126 394572 397132 394574
rect 397196 394572 397202 394636
rect 217726 393892 217732 393956
rect 217796 393954 217802 393956
rect 218145 393954 218211 393957
rect 217796 393952 218211 393954
rect 217796 393896 218150 393952
rect 218206 393896 218211 393952
rect 217796 393894 218211 393896
rect 217796 393892 217802 393894
rect 218145 393891 218211 393894
rect 39021 393546 39087 393549
rect 39990 393546 40050 393766
rect 217174 393756 217180 393820
rect 217244 393818 217250 393820
rect 218605 393818 218671 393821
rect 396625 393818 396691 393821
rect 217244 393816 219450 393818
rect 217244 393760 218610 393816
rect 218666 393796 219450 393816
rect 396625 393816 399402 393818
rect 218666 393760 220064 393796
rect 217244 393758 220064 393760
rect 217244 393756 217250 393758
rect 218605 393755 218671 393758
rect 219390 393736 220064 393758
rect 396625 393760 396630 393816
rect 396686 393796 399402 393816
rect 396686 393760 400016 393796
rect 396625 393758 400016 393760
rect 396625 393755 396691 393758
rect 399342 393736 400016 393758
rect 39021 393544 40050 393546
rect 39021 393488 39026 393544
rect 39082 393488 40050 393544
rect 39021 393486 40050 393488
rect 39021 393483 39087 393486
rect 217133 392866 217199 392869
rect 218513 392866 218579 392869
rect 396993 392866 397059 392869
rect 217133 392864 219450 392866
rect 38837 392322 38903 392325
rect 39990 392322 40050 392814
rect 217133 392808 217138 392864
rect 217194 392808 218518 392864
rect 218574 392844 219450 392864
rect 396993 392864 399402 392866
rect 218574 392808 220064 392844
rect 217133 392806 220064 392808
rect 217133 392803 217199 392806
rect 218513 392803 218579 392806
rect 219390 392784 220064 392806
rect 396993 392808 396998 392864
rect 397054 392844 399402 392864
rect 397054 392808 400016 392844
rect 396993 392806 400016 392808
rect 396993 392803 397059 392806
rect 399342 392784 400016 392806
rect 38837 392320 40050 392322
rect 38837 392264 38842 392320
rect 38898 392264 40050 392320
rect 38837 392262 40050 392264
rect 38837 392259 38903 392262
rect 216949 391914 217015 391917
rect 217225 391914 217291 391917
rect 216949 391912 217291 391914
rect 216949 391856 216954 391912
rect 217010 391856 217230 391912
rect 217286 391856 217291 391912
rect 216949 391854 217291 391856
rect 216949 391851 217015 391854
rect 217225 391851 217291 391854
rect 583520 391628 584960 391868
rect 216949 391098 217015 391101
rect 397085 391098 397151 391101
rect 216949 391096 219450 391098
rect 38929 390690 38995 390693
rect 39990 390690 40050 391046
rect 216949 391040 216954 391096
rect 217010 391076 219450 391096
rect 397085 391096 399402 391098
rect 217010 391040 220064 391076
rect 216949 391038 220064 391040
rect 216949 391035 217015 391038
rect 219390 391016 220064 391038
rect 397085 391040 397090 391096
rect 397146 391076 399402 391096
rect 397146 391040 400016 391076
rect 397085 391038 400016 391040
rect 397085 391035 397151 391038
rect 399342 391016 400016 391038
rect 38929 390688 40050 390690
rect 38929 390632 38934 390688
rect 38990 390632 40050 390688
rect 38929 390630 40050 390632
rect 38929 390627 38995 390630
rect 216857 390554 216923 390557
rect 217869 390554 217935 390557
rect 216857 390552 217935 390554
rect 216857 390496 216862 390552
rect 216918 390496 217874 390552
rect 217930 390496 217935 390552
rect 216857 390494 217935 390496
rect 216857 390491 216923 390494
rect 217869 390491 217935 390494
rect 217869 390010 217935 390013
rect 396901 390010 396967 390013
rect 217869 390008 219450 390010
rect 38745 389466 38811 389469
rect 39990 389466 40050 389958
rect 217869 389952 217874 390008
rect 217930 389988 219450 390008
rect 396901 390008 399402 390010
rect 217930 389952 220064 389988
rect 217869 389950 220064 389952
rect 217869 389947 217935 389950
rect 219390 389928 220064 389950
rect 396901 389952 396906 390008
rect 396962 389988 399402 390008
rect 396962 389952 400016 389988
rect 396901 389950 400016 389952
rect 396901 389947 396967 389950
rect 399342 389928 400016 389950
rect 38745 389464 40050 389466
rect 38745 389408 38750 389464
rect 38806 389408 40050 389464
rect 38745 389406 40050 389408
rect 38745 389403 38811 389406
rect 217225 388242 217291 388245
rect 217409 388242 217475 388245
rect 396809 388242 396875 388245
rect 217225 388240 219450 388242
rect 38653 387834 38719 387837
rect 39990 387834 40050 388190
rect 217225 388184 217230 388240
rect 217286 388184 217414 388240
rect 217470 388220 219450 388240
rect 396809 388240 399402 388242
rect 217470 388184 220064 388220
rect 217225 388182 220064 388184
rect 217225 388179 217291 388182
rect 217409 388179 217475 388182
rect 219390 388160 220064 388182
rect 396809 388184 396814 388240
rect 396870 388220 399402 388240
rect 396870 388184 400016 388220
rect 396809 388182 400016 388184
rect 396809 388179 396875 388182
rect 399342 388160 400016 388182
rect 38653 387832 40050 387834
rect 38653 387776 38658 387832
rect 38714 387776 40050 387832
rect 38653 387774 40050 387776
rect 38653 387771 38719 387774
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 216673 370018 216739 370021
rect 217358 370018 217364 370020
rect 216673 370016 217364 370018
rect 38561 369882 38627 369885
rect 39990 369882 40050 369966
rect 216673 369960 216678 370016
rect 216734 369960 217364 370016
rect 216673 369958 217364 369960
rect 216673 369955 216739 369958
rect 217358 369956 217364 369958
rect 217428 370018 217434 370020
rect 396441 370018 396507 370021
rect 396717 370018 396783 370021
rect 217428 369996 219450 370018
rect 396441 370016 399402 370018
rect 217428 369958 220064 369996
rect 217428 369956 217434 369958
rect 219390 369936 220064 369958
rect 396441 369960 396446 370016
rect 396502 369960 396722 370016
rect 396778 369996 399402 370016
rect 396778 369960 400016 369996
rect 396441 369958 400016 369960
rect 396441 369955 396507 369958
rect 396717 369955 396783 369958
rect 399342 369936 400016 369958
rect 216857 369884 216923 369885
rect 216806 369882 216812 369884
rect 38561 369880 40050 369882
rect 38561 369824 38566 369880
rect 38622 369824 40050 369880
rect 38561 369822 40050 369824
rect 216766 369822 216812 369882
rect 216876 369880 216923 369884
rect 216918 369824 216923 369880
rect 38561 369819 38627 369822
rect 216806 369820 216812 369822
rect 216876 369820 216923 369824
rect 216857 369819 216923 369820
rect 37733 368386 37799 368389
rect 38193 368386 38259 368389
rect 216857 368386 216923 368389
rect 217542 368386 217548 368388
rect 37733 368384 40050 368386
rect 37733 368328 37738 368384
rect 37794 368328 38198 368384
rect 38254 368328 40050 368384
rect 37733 368326 40050 368328
rect 216857 368384 217548 368386
rect 216857 368328 216862 368384
rect 216918 368328 217548 368384
rect 216857 368326 217548 368328
rect 37733 368323 37799 368326
rect 38193 368323 38259 368326
rect 216857 368323 216923 368326
rect 217542 368324 217548 368326
rect 217612 368324 217618 368388
rect 217910 368324 217916 368388
rect 217980 368386 217986 368388
rect 218513 368386 218579 368389
rect 396717 368386 396783 368389
rect 397310 368386 397316 368388
rect 217980 368384 219450 368386
rect 217980 368328 218518 368384
rect 218574 368364 219450 368384
rect 396717 368384 397316 368386
rect 218574 368328 220064 368364
rect 217980 368326 220064 368328
rect 217980 368324 217986 368326
rect 218513 368323 218579 368326
rect 219390 368304 220064 368326
rect 396717 368328 396722 368384
rect 396778 368328 397316 368384
rect 396717 368326 397316 368328
rect 396717 368323 396783 368326
rect 397310 368324 397316 368326
rect 397380 368386 397386 368388
rect 397380 368364 399402 368386
rect 397380 368326 400016 368364
rect 397380 368324 397386 368326
rect 399342 368304 400016 368326
rect 217409 368114 217475 368117
rect 396533 368114 396599 368117
rect 217409 368112 219450 368114
rect 38377 367570 38443 367573
rect 39990 367570 40050 368062
rect 217409 368056 217414 368112
rect 217470 368092 219450 368112
rect 396533 368112 399402 368114
rect 217470 368056 220064 368092
rect 217409 368054 220064 368056
rect 217409 368051 217475 368054
rect 219390 368032 220064 368054
rect 396533 368056 396538 368112
rect 396594 368092 399402 368112
rect 396594 368056 400016 368092
rect 396533 368054 400016 368056
rect 396533 368051 396599 368054
rect 399342 368032 400016 368054
rect 38377 367568 40050 367570
rect 38377 367512 38382 367568
rect 38438 367512 40050 367568
rect 38377 367510 40050 367512
rect 38377 367507 38443 367510
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect 219198 359892 219204 359956
rect 219268 359954 219274 359956
rect 221917 359954 221983 359957
rect 219268 359952 221983 359954
rect 219268 359896 221922 359952
rect 221978 359896 221983 359952
rect 219268 359894 221983 359896
rect 219268 359892 219274 359894
rect 221917 359891 221983 359894
rect 217726 359620 217732 359684
rect 217796 359682 217802 359684
rect 263869 359682 263935 359685
rect 217796 359680 263935 359682
rect 217796 359624 263874 359680
rect 263930 359624 263935 359680
rect 217796 359622 263935 359624
rect 217796 359620 217802 359622
rect 263869 359619 263935 359622
rect 212349 359546 212415 359549
rect 253197 359546 253263 359549
rect 212349 359544 253263 359546
rect 212349 359488 212354 359544
rect 212410 359488 253202 359544
rect 253258 359488 253263 359544
rect 212349 359486 253263 359488
rect 212349 359483 212415 359486
rect 253197 359483 253263 359486
rect 285213 359546 285279 359549
rect 357566 359546 357572 359548
rect 285213 359544 357572 359546
rect 285213 359488 285218 359544
rect 285274 359488 357572 359544
rect 285213 359486 357572 359488
rect 285213 359483 285279 359486
rect 357566 359484 357572 359486
rect 357636 359484 357642 359548
rect 450854 359484 450860 359548
rect 450924 359546 450930 359548
rect 451136 359546 451142 359548
rect 450924 359486 451142 359546
rect 450924 359484 450930 359486
rect 451136 359484 451142 359486
rect 451206 359484 451212 359548
rect 218830 359348 218836 359412
rect 218900 359410 218906 359412
rect 266629 359410 266695 359413
rect 218900 359408 266695 359410
rect 218900 359352 266634 359408
rect 266690 359352 266695 359408
rect 218900 359350 266695 359352
rect 218900 359348 218906 359350
rect 266629 359347 266695 359350
rect 282269 359410 282335 359413
rect 358854 359410 358860 359412
rect 282269 359408 358860 359410
rect 282269 359352 282274 359408
rect 282330 359352 358860 359408
rect 282269 359350 358860 359352
rect 282269 359347 282335 359350
rect 358854 359348 358860 359350
rect 358924 359348 358930 359412
rect 253197 359274 253263 359277
rect 260557 359274 260623 359277
rect 253197 359272 260623 359274
rect 253197 359216 253202 359272
rect 253258 359216 260562 359272
rect 260618 359216 260623 359272
rect 253197 359214 260623 359216
rect 253197 359211 253263 359214
rect 260557 359211 260623 359214
rect 216254 358668 216260 358732
rect 216324 358730 216330 358732
rect 223757 358730 223823 358733
rect 216324 358728 223823 358730
rect 216324 358672 223762 358728
rect 223818 358672 223823 358728
rect 216324 358670 223823 358672
rect 216324 358668 216330 358670
rect 223757 358667 223823 358670
rect 325693 358730 325759 358733
rect 325918 358730 325924 358732
rect 325693 358728 325924 358730
rect 325693 358672 325698 358728
rect 325754 358672 325924 358728
rect 325693 358670 325924 358672
rect 325693 358667 325759 358670
rect 325918 358668 325924 358670
rect 325988 358668 325994 358732
rect 216581 358594 216647 358597
rect 228173 358594 228239 358597
rect 235993 358596 236059 358597
rect 235942 358594 235948 358596
rect 216581 358592 228239 358594
rect -960 358458 480 358548
rect 216581 358536 216586 358592
rect 216642 358536 228178 358592
rect 228234 358536 228239 358592
rect 216581 358534 228239 358536
rect 235902 358534 235948 358594
rect 236012 358592 236059 358596
rect 236054 358536 236059 358592
rect 216581 358531 216647 358534
rect 228173 358531 228239 358534
rect 235942 358532 235948 358534
rect 236012 358532 236059 358536
rect 235993 358531 236059 358532
rect 308765 358594 308831 358597
rect 359089 358594 359155 358597
rect 308765 358592 359155 358594
rect 308765 358536 308770 358592
rect 308826 358536 359094 358592
rect 359150 358536 359155 358592
rect 308765 358534 359155 358536
rect 308765 358531 308831 358534
rect 359089 358531 359155 358534
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 210734 358396 210740 358460
rect 210804 358458 210810 358460
rect 219341 358458 219407 358461
rect 210804 358456 219407 358458
rect 210804 358400 219346 358456
rect 219402 358400 219407 358456
rect 210804 358398 219407 358400
rect 210804 358396 210810 358398
rect 219341 358395 219407 358398
rect 224217 358458 224283 358461
rect 234061 358458 234127 358461
rect 224217 358456 234127 358458
rect 224217 358400 224222 358456
rect 224278 358400 234066 358456
rect 234122 358400 234127 358456
rect 224217 358398 234127 358400
rect 224217 358395 224283 358398
rect 234061 358395 234127 358398
rect 305821 358458 305887 358461
rect 357709 358458 357775 358461
rect 305821 358456 357775 358458
rect 305821 358400 305826 358456
rect 305882 358400 357714 358456
rect 357770 358400 357775 358456
rect 305821 358398 357775 358400
rect 305821 358395 305887 358398
rect 357709 358395 357775 358398
rect 213545 358322 213611 358325
rect 232221 358322 232287 358325
rect 213545 358320 232287 358322
rect 213545 358264 213550 358320
rect 213606 358264 232226 358320
rect 232282 358264 232287 358320
rect 213545 358262 232287 358264
rect 213545 358259 213611 358262
rect 232221 358259 232287 358262
rect 299933 358322 299999 358325
rect 357525 358322 357591 358325
rect 299933 358320 357591 358322
rect 299933 358264 299938 358320
rect 299994 358264 357530 358320
rect 357586 358264 357591 358320
rect 299933 358262 357591 358264
rect 299933 358259 299999 358262
rect 357525 358259 357591 358262
rect 60590 358124 60596 358188
rect 60660 358186 60666 358188
rect 61377 358186 61443 358189
rect 64321 358188 64387 358189
rect 60660 358184 61443 358186
rect 60660 358128 61382 358184
rect 61438 358128 61443 358184
rect 60660 358126 61443 358128
rect 60660 358124 60666 358126
rect 61377 358123 61443 358126
rect 64270 358124 64276 358188
rect 64340 358186 64387 358188
rect 64340 358184 64432 358186
rect 64382 358128 64432 358184
rect 64340 358126 64432 358128
rect 64340 358124 64387 358126
rect 219014 358124 219020 358188
rect 219084 358186 219090 358188
rect 250621 358186 250687 358189
rect 276013 358188 276079 358189
rect 300853 358188 300919 358189
rect 276013 358186 276060 358188
rect 219084 358184 250687 358186
rect 219084 358128 250626 358184
rect 250682 358128 250687 358184
rect 219084 358126 250687 358128
rect 275968 358184 276060 358186
rect 275968 358128 276018 358184
rect 275968 358126 276060 358128
rect 219084 358124 219090 358126
rect 64321 358123 64387 358124
rect 250621 358123 250687 358126
rect 276013 358124 276060 358126
rect 276124 358124 276130 358188
rect 300853 358186 300900 358188
rect 300808 358184 300900 358186
rect 300808 358128 300858 358184
rect 300808 358126 300900 358128
rect 300853 358124 300900 358126
rect 300964 358124 300970 358188
rect 301037 358186 301103 358189
rect 357617 358186 357683 358189
rect 416037 358188 416103 358189
rect 488533 358188 488599 358189
rect 416037 358186 416084 358188
rect 301037 358184 357683 358186
rect 301037 358128 301042 358184
rect 301098 358128 357622 358184
rect 357678 358128 357683 358184
rect 301037 358126 357683 358128
rect 415992 358184 416084 358186
rect 415992 358128 416042 358184
rect 415992 358126 416084 358128
rect 276013 358123 276079 358124
rect 300853 358123 300919 358124
rect 301037 358123 301103 358126
rect 357617 358123 357683 358126
rect 416037 358124 416084 358126
rect 416148 358124 416154 358188
rect 488533 358186 488580 358188
rect 488488 358184 488580 358186
rect 488488 358128 488538 358184
rect 488488 358126 488580 358128
rect 488533 358124 488580 358126
rect 488644 358124 488650 358188
rect 416037 358123 416103 358124
rect 488533 358123 488599 358124
rect 219985 358050 220051 358053
rect 253933 358050 253999 358053
rect 219985 358048 253999 358050
rect 219985 357992 219990 358048
rect 220046 357992 253938 358048
rect 253994 357992 253999 358048
rect 219985 357990 253999 357992
rect 219985 357987 220051 357990
rect 253933 357987 253999 357990
rect 294045 358050 294111 358053
rect 356605 358050 356671 358053
rect 294045 358048 356671 358050
rect 294045 357992 294050 358048
rect 294106 357992 356610 358048
rect 356666 357992 356671 358048
rect 294045 357990 356671 357992
rect 294045 357987 294111 357990
rect 356605 357987 356671 357990
rect 296989 357914 297055 357917
rect 301037 357914 301103 357917
rect 296989 357912 301103 357914
rect 296989 357856 296994 357912
rect 297050 357856 301042 357912
rect 301098 357856 301103 357912
rect 296989 357854 301103 357856
rect 296989 357851 297055 357854
rect 301037 357851 301103 357854
rect 55990 357308 55996 357372
rect 56060 357370 56066 357372
rect 56501 357370 56567 357373
rect 56060 357368 56567 357370
rect 56060 357312 56506 357368
rect 56562 357312 56567 357368
rect 56060 357310 56567 357312
rect 56060 357308 56066 357310
rect 56501 357307 56567 357310
rect 58198 357308 58204 357372
rect 58268 357370 58274 357372
rect 59261 357370 59327 357373
rect 58268 357368 59327 357370
rect 58268 357312 59266 357368
rect 59322 357312 59327 357368
rect 58268 357310 59327 357312
rect 58268 357308 58274 357310
rect 59261 357307 59327 357310
rect 59670 357308 59676 357372
rect 59740 357370 59746 357372
rect 60641 357370 60707 357373
rect 59740 357368 60707 357370
rect 59740 357312 60646 357368
rect 60702 357312 60707 357368
rect 59740 357310 60707 357312
rect 59740 357308 59746 357310
rect 60641 357307 60707 357310
rect 61878 357308 61884 357372
rect 61948 357370 61954 357372
rect 62021 357370 62087 357373
rect 61948 357368 62087 357370
rect 61948 357312 62026 357368
rect 62082 357312 62087 357368
rect 61948 357310 62087 357312
rect 61948 357308 61954 357310
rect 62021 357307 62087 357310
rect 63166 357308 63172 357372
rect 63236 357370 63242 357372
rect 63401 357370 63467 357373
rect 63236 357368 63467 357370
rect 63236 357312 63406 357368
rect 63462 357312 63467 357368
rect 63236 357310 63467 357312
rect 63236 357308 63242 357310
rect 63401 357307 63467 357310
rect 66478 357308 66484 357372
rect 66548 357370 66554 357372
rect 67541 357370 67607 357373
rect 66548 357368 67607 357370
rect 66548 357312 67546 357368
rect 67602 357312 67607 357368
rect 66548 357310 67607 357312
rect 66548 357308 66554 357310
rect 67541 357307 67607 357310
rect 68686 357308 68692 357372
rect 68756 357370 68762 357372
rect 68829 357370 68895 357373
rect 68756 357368 68895 357370
rect 68756 357312 68834 357368
rect 68890 357312 68895 357368
rect 68756 357310 68895 357312
rect 68756 357308 68762 357310
rect 68829 357307 68895 357310
rect 70158 357308 70164 357372
rect 70228 357370 70234 357372
rect 70301 357370 70367 357373
rect 70228 357368 70367 357370
rect 70228 357312 70306 357368
rect 70362 357312 70367 357368
rect 70228 357310 70367 357312
rect 70228 357308 70234 357310
rect 70301 357307 70367 357310
rect 71262 357308 71268 357372
rect 71332 357370 71338 357372
rect 71681 357370 71747 357373
rect 71332 357368 71747 357370
rect 71332 357312 71686 357368
rect 71742 357312 71747 357368
rect 71332 357310 71747 357312
rect 71332 357308 71338 357310
rect 71681 357307 71747 357310
rect 72366 357308 72372 357372
rect 72436 357370 72442 357372
rect 73061 357370 73127 357373
rect 72436 357368 73127 357370
rect 72436 357312 73066 357368
rect 73122 357312 73127 357368
rect 72436 357310 73127 357312
rect 72436 357308 72442 357310
rect 73061 357307 73127 357310
rect 73470 357308 73476 357372
rect 73540 357370 73546 357372
rect 74349 357370 74415 357373
rect 73540 357368 74415 357370
rect 73540 357312 74354 357368
rect 74410 357312 74415 357368
rect 73540 357310 74415 357312
rect 73540 357308 73546 357310
rect 74349 357307 74415 357310
rect 74574 357308 74580 357372
rect 74644 357370 74650 357372
rect 75821 357370 75887 357373
rect 74644 357368 75887 357370
rect 74644 357312 75826 357368
rect 75882 357312 75887 357368
rect 74644 357310 75887 357312
rect 74644 357308 74650 357310
rect 75821 357307 75887 357310
rect 76005 357370 76071 357373
rect 76966 357370 76972 357372
rect 76005 357368 76972 357370
rect 76005 357312 76010 357368
rect 76066 357312 76972 357368
rect 76005 357310 76972 357312
rect 76005 357307 76071 357310
rect 76966 357308 76972 357310
rect 77036 357308 77042 357372
rect 78438 357308 78444 357372
rect 78508 357370 78514 357372
rect 78581 357370 78647 357373
rect 78508 357368 78647 357370
rect 78508 357312 78586 357368
rect 78642 357312 78647 357368
rect 78508 357310 78647 357312
rect 78508 357308 78514 357310
rect 78581 357307 78647 357310
rect 79542 357308 79548 357372
rect 79612 357370 79618 357372
rect 79961 357370 80027 357373
rect 79612 357368 80027 357370
rect 79612 357312 79966 357368
rect 80022 357312 80027 357368
rect 79612 357310 80027 357312
rect 79612 357308 79618 357310
rect 79961 357307 80027 357310
rect 81014 357308 81020 357372
rect 81084 357370 81090 357372
rect 81341 357370 81407 357373
rect 81084 357368 81407 357370
rect 81084 357312 81346 357368
rect 81402 357312 81407 357368
rect 81084 357310 81407 357312
rect 81084 357308 81090 357310
rect 81341 357307 81407 357310
rect 85982 357308 85988 357372
rect 86052 357370 86058 357372
rect 86861 357370 86927 357373
rect 88241 357372 88307 357373
rect 91001 357372 91067 357373
rect 86052 357368 86927 357370
rect 86052 357312 86866 357368
rect 86922 357312 86927 357368
rect 86052 357310 86927 357312
rect 86052 357308 86058 357310
rect 86861 357307 86927 357310
rect 88190 357308 88196 357372
rect 88260 357370 88307 357372
rect 88260 357368 88352 357370
rect 88302 357312 88352 357368
rect 88260 357310 88352 357312
rect 88260 357308 88307 357310
rect 90950 357308 90956 357372
rect 91020 357370 91067 357372
rect 93393 357370 93459 357373
rect 93526 357370 93532 357372
rect 91020 357368 91112 357370
rect 91062 357312 91112 357368
rect 91020 357310 91112 357312
rect 93393 357368 93532 357370
rect 93393 357312 93398 357368
rect 93454 357312 93532 357368
rect 93393 357310 93532 357312
rect 91020 357308 91067 357310
rect 88241 357307 88307 357308
rect 91001 357307 91067 357308
rect 93393 357307 93459 357310
rect 93526 357308 93532 357310
rect 93596 357308 93602 357372
rect 95918 357308 95924 357372
rect 95988 357370 95994 357372
rect 96521 357370 96587 357373
rect 95988 357368 96587 357370
rect 95988 357312 96526 357368
rect 96582 357312 96587 357368
rect 95988 357310 96587 357312
rect 95988 357308 95994 357310
rect 96521 357307 96587 357310
rect 98494 357308 98500 357372
rect 98564 357370 98570 357372
rect 99281 357370 99347 357373
rect 98564 357368 99347 357370
rect 98564 357312 99286 357368
rect 99342 357312 99347 357368
rect 98564 357310 99347 357312
rect 98564 357308 98570 357310
rect 99281 357307 99347 357310
rect 100886 357308 100892 357372
rect 100956 357370 100962 357372
rect 102041 357370 102107 357373
rect 100956 357368 102107 357370
rect 100956 357312 102046 357368
rect 102102 357312 102107 357368
rect 100956 357310 102107 357312
rect 100956 357308 100962 357310
rect 102041 357307 102107 357310
rect 106038 357308 106044 357372
rect 106108 357370 106114 357372
rect 106181 357370 106247 357373
rect 106108 357368 106247 357370
rect 106108 357312 106186 357368
rect 106242 357312 106247 357368
rect 106108 357310 106247 357312
rect 106108 357308 106114 357310
rect 106181 357307 106247 357310
rect 243118 357308 243124 357372
rect 243188 357370 243194 357372
rect 243537 357370 243603 357373
rect 243188 357368 243603 357370
rect 243188 357312 243542 357368
rect 243598 357312 243603 357368
rect 243188 357310 243603 357312
rect 243188 357308 243194 357310
rect 243537 357307 243603 357310
rect 247217 357370 247283 357373
rect 248689 357372 248755 357373
rect 248270 357370 248276 357372
rect 247217 357368 248276 357370
rect 247217 357312 247222 357368
rect 247278 357312 248276 357368
rect 247217 357310 248276 357312
rect 247217 357307 247283 357310
rect 248270 357308 248276 357310
rect 248340 357308 248346 357372
rect 248638 357370 248644 357372
rect 248598 357310 248644 357370
rect 248708 357368 248755 357372
rect 248750 357312 248755 357368
rect 248638 357308 248644 357310
rect 248708 357308 248755 357312
rect 248689 357307 248755 357308
rect 249977 357370 250043 357373
rect 251265 357372 251331 357373
rect 250662 357370 250668 357372
rect 249977 357368 250668 357370
rect 249977 357312 249982 357368
rect 250038 357312 250668 357368
rect 249977 357310 250668 357312
rect 249977 357307 250043 357310
rect 250662 357308 250668 357310
rect 250732 357308 250738 357372
rect 251214 357370 251220 357372
rect 251174 357310 251220 357370
rect 251284 357368 251331 357372
rect 251326 357312 251331 357368
rect 251214 357308 251220 357310
rect 251284 357308 251331 357312
rect 251265 357307 251331 357308
rect 252645 357370 252711 357373
rect 254577 357372 254643 357373
rect 253606 357370 253612 357372
rect 252645 357368 253612 357370
rect 252645 357312 252650 357368
rect 252706 357312 253612 357368
rect 252645 357310 253612 357312
rect 252645 357307 252711 357310
rect 253606 357308 253612 357310
rect 253676 357308 253682 357372
rect 254526 357370 254532 357372
rect 254486 357310 254532 357370
rect 254596 357368 254643 357372
rect 254638 357312 254643 357368
rect 254526 357308 254532 357310
rect 254596 357308 254643 357312
rect 254577 357307 254643 357308
rect 255405 357370 255471 357373
rect 255998 357370 256004 357372
rect 255405 357368 256004 357370
rect 255405 357312 255410 357368
rect 255466 357312 256004 357368
rect 255405 357310 256004 357312
rect 255405 357307 255471 357310
rect 255998 357308 256004 357310
rect 256068 357308 256074 357372
rect 257102 357308 257108 357372
rect 257172 357370 257178 357372
rect 257337 357370 257403 357373
rect 257172 357368 257403 357370
rect 257172 357312 257342 357368
rect 257398 357312 257403 357368
rect 257172 357310 257403 357312
rect 257172 357308 257178 357310
rect 257337 357307 257403 357310
rect 258165 357370 258231 357373
rect 258390 357370 258396 357372
rect 258165 357368 258396 357370
rect 258165 357312 258170 357368
rect 258226 357312 258396 357368
rect 258165 357310 258396 357312
rect 258165 357307 258231 357310
rect 258390 357308 258396 357310
rect 258460 357308 258466 357372
rect 260833 357370 260899 357373
rect 262121 357372 262187 357373
rect 260966 357370 260972 357372
rect 260833 357368 260972 357370
rect 260833 357312 260838 357368
rect 260894 357312 260972 357368
rect 260833 357310 260972 357312
rect 260833 357307 260899 357310
rect 260966 357308 260972 357310
rect 261036 357308 261042 357372
rect 262070 357370 262076 357372
rect 262030 357310 262076 357370
rect 262140 357368 262187 357372
rect 262182 357312 262187 357368
rect 262070 357308 262076 357310
rect 262140 357308 262187 357312
rect 262121 357307 262187 357308
rect 262765 357372 262831 357373
rect 262765 357368 262812 357372
rect 262876 357370 262882 357372
rect 262765 357312 262770 357368
rect 262765 357308 262812 357312
rect 262876 357310 262922 357370
rect 262876 357308 262882 357310
rect 263542 357308 263548 357372
rect 263612 357370 263618 357372
rect 263685 357370 263751 357373
rect 263961 357372 264027 357373
rect 263612 357368 263751 357370
rect 263612 357312 263690 357368
rect 263746 357312 263751 357368
rect 263612 357310 263751 357312
rect 263612 357308 263618 357310
rect 262765 357307 262831 357308
rect 263685 357307 263751 357310
rect 263910 357308 263916 357372
rect 263980 357370 264027 357372
rect 265709 357372 265775 357373
rect 263980 357368 264072 357370
rect 264022 357312 264072 357368
rect 263980 357310 264072 357312
rect 265709 357368 265756 357372
rect 265820 357370 265826 357372
rect 265709 357312 265714 357368
rect 263980 357308 264027 357310
rect 263961 357307 264027 357308
rect 265709 357308 265756 357312
rect 265820 357310 265866 357370
rect 265820 357308 265826 357310
rect 266302 357308 266308 357372
rect 266372 357370 266378 357372
rect 266445 357370 266511 357373
rect 267549 357372 267615 357373
rect 267549 357370 267596 357372
rect 266372 357368 266511 357370
rect 266372 357312 266450 357368
rect 266506 357312 266511 357368
rect 266372 357310 266511 357312
rect 267504 357368 267596 357370
rect 267504 357312 267554 357368
rect 267504 357310 267596 357312
rect 266372 357308 266378 357310
rect 265709 357307 265775 357308
rect 266445 357307 266511 357310
rect 267549 357308 267596 357310
rect 267660 357308 267666 357372
rect 267733 357370 267799 357373
rect 268561 357372 268627 357373
rect 268326 357370 268332 357372
rect 267733 357368 268332 357370
rect 267733 357312 267738 357368
rect 267794 357312 268332 357368
rect 267733 357310 268332 357312
rect 267549 357307 267615 357308
rect 267733 357307 267799 357310
rect 268326 357308 268332 357310
rect 268396 357308 268402 357372
rect 268510 357308 268516 357372
rect 268580 357370 268627 357372
rect 269757 357372 269823 357373
rect 268580 357368 268672 357370
rect 268622 357312 268672 357368
rect 268580 357310 268672 357312
rect 269757 357368 269804 357372
rect 269868 357370 269874 357372
rect 270585 357370 270651 357373
rect 271137 357372 271203 357373
rect 270902 357370 270908 357372
rect 269757 357312 269762 357368
rect 268580 357308 268627 357310
rect 268561 357307 268627 357308
rect 269757 357308 269804 357312
rect 269868 357310 269914 357370
rect 270585 357368 270908 357370
rect 270585 357312 270590 357368
rect 270646 357312 270908 357368
rect 270585 357310 270908 357312
rect 269868 357308 269874 357310
rect 269757 357307 269823 357308
rect 270585 357307 270651 357310
rect 270902 357308 270908 357310
rect 270972 357308 270978 357372
rect 271086 357308 271092 357372
rect 271156 357370 271203 357372
rect 272149 357372 272215 357373
rect 273345 357372 273411 357373
rect 271156 357368 271248 357370
rect 271198 357312 271248 357368
rect 271156 357310 271248 357312
rect 272149 357368 272196 357372
rect 272260 357370 272266 357372
rect 273294 357370 273300 357372
rect 272149 357312 272154 357368
rect 271156 357308 271203 357310
rect 271137 357307 271203 357308
rect 272149 357308 272196 357312
rect 272260 357310 272306 357370
rect 273254 357310 273300 357370
rect 273364 357368 273411 357372
rect 273406 357312 273411 357368
rect 272260 357308 272266 357310
rect 273294 357308 273300 357310
rect 273364 357308 273411 357312
rect 274398 357308 274404 357372
rect 274468 357370 274474 357372
rect 274541 357370 274607 357373
rect 275921 357372 275987 357373
rect 277025 357372 277091 357373
rect 275870 357370 275876 357372
rect 274468 357368 274607 357370
rect 274468 357312 274546 357368
rect 274602 357312 274607 357368
rect 274468 357310 274607 357312
rect 275830 357310 275876 357370
rect 275940 357368 275987 357372
rect 276974 357370 276980 357372
rect 275982 357312 275987 357368
rect 274468 357308 274474 357310
rect 272149 357307 272215 357308
rect 273345 357307 273411 357308
rect 274541 357307 274607 357310
rect 275870 357308 275876 357310
rect 275940 357308 275987 357312
rect 276934 357310 276980 357370
rect 277044 357368 277091 357372
rect 277086 357312 277091 357368
rect 276974 357308 276980 357310
rect 277044 357308 277091 357312
rect 275921 357307 275987 357308
rect 277025 357307 277091 357308
rect 282913 357370 282979 357373
rect 283414 357370 283420 357372
rect 282913 357368 283420 357370
rect 282913 357312 282918 357368
rect 282974 357312 283420 357368
rect 282913 357310 283420 357312
rect 282913 357307 282979 357310
rect 283414 357308 283420 357310
rect 283484 357308 283490 357372
rect 285673 357370 285739 357373
rect 285990 357370 285996 357372
rect 285673 357368 285996 357370
rect 285673 357312 285678 357368
rect 285734 357312 285996 357368
rect 285673 357310 285996 357312
rect 285673 357307 285739 357310
rect 285990 357308 285996 357310
rect 286060 357308 286066 357372
rect 287053 357370 287119 357373
rect 288198 357370 288204 357372
rect 287053 357368 288204 357370
rect 287053 357312 287058 357368
rect 287114 357312 288204 357368
rect 287053 357310 288204 357312
rect 287053 357307 287119 357310
rect 288198 357308 288204 357310
rect 288268 357308 288274 357372
rect 289905 357370 289971 357373
rect 290958 357370 290964 357372
rect 289905 357368 290964 357370
rect 289905 357312 289910 357368
rect 289966 357312 290964 357368
rect 289905 357310 290964 357312
rect 289905 357307 289971 357310
rect 290958 357308 290964 357310
rect 291028 357308 291034 357372
rect 292573 357370 292639 357373
rect 293350 357370 293356 357372
rect 292573 357368 293356 357370
rect 292573 357312 292578 357368
rect 292634 357312 293356 357368
rect 292573 357310 293356 357312
rect 292573 357307 292639 357310
rect 293350 357308 293356 357310
rect 293420 357308 293426 357372
rect 295333 357370 295399 357373
rect 295926 357370 295932 357372
rect 295333 357368 295932 357370
rect 295333 357312 295338 357368
rect 295394 357312 295932 357368
rect 295333 357310 295932 357312
rect 295333 357307 295399 357310
rect 295926 357308 295932 357310
rect 295996 357308 296002 357372
rect 298185 357370 298251 357373
rect 298502 357370 298508 357372
rect 298185 357368 298508 357370
rect 298185 357312 298190 357368
rect 298246 357312 298508 357368
rect 298185 357310 298508 357312
rect 298185 357307 298251 357310
rect 298502 357308 298508 357310
rect 298572 357308 298578 357372
rect 302233 357370 302299 357373
rect 303470 357370 303476 357372
rect 302233 357368 303476 357370
rect 302233 357312 302238 357368
rect 302294 357312 303476 357368
rect 302233 357310 303476 357312
rect 302233 357307 302299 357310
rect 303470 357308 303476 357310
rect 303540 357308 303546 357372
rect 304993 357370 305059 357373
rect 305862 357370 305868 357372
rect 304993 357368 305868 357370
rect 304993 357312 304998 357368
rect 305054 357312 305868 357368
rect 304993 357310 305868 357312
rect 304993 357307 305059 357310
rect 305862 357308 305868 357310
rect 305932 357308 305938 357372
rect 307753 357370 307819 357373
rect 308070 357370 308076 357372
rect 307753 357368 308076 357370
rect 307753 357312 307758 357368
rect 307814 357312 308076 357368
rect 307753 357310 308076 357312
rect 307753 357307 307819 357310
rect 308070 357308 308076 357310
rect 308140 357308 308146 357372
rect 310513 357370 310579 357373
rect 311014 357370 311020 357372
rect 310513 357368 311020 357370
rect 310513 357312 310518 357368
rect 310574 357312 311020 357368
rect 310513 357310 311020 357312
rect 310513 357307 310579 357310
rect 311014 357308 311020 357310
rect 311084 357308 311090 357372
rect 313273 357370 313339 357373
rect 313406 357370 313412 357372
rect 313273 357368 313412 357370
rect 313273 357312 313278 357368
rect 313334 357312 313412 357368
rect 313273 357310 313412 357312
rect 313273 357307 313339 357310
rect 313406 357308 313412 357310
rect 313476 357308 313482 357372
rect 314745 357370 314811 357373
rect 315614 357370 315620 357372
rect 314745 357368 315620 357370
rect 314745 357312 314750 357368
rect 314806 357312 315620 357368
rect 314745 357310 315620 357312
rect 314745 357307 314811 357310
rect 315614 357308 315620 357310
rect 315684 357308 315690 357372
rect 317413 357370 317479 357373
rect 318374 357370 318380 357372
rect 317413 357368 318380 357370
rect 317413 357312 317418 357368
rect 317474 357312 318380 357368
rect 317413 357310 318380 357312
rect 317413 357307 317479 357310
rect 318374 357308 318380 357310
rect 318444 357308 318450 357372
rect 320173 357370 320239 357373
rect 320950 357370 320956 357372
rect 320173 357368 320956 357370
rect 320173 357312 320178 357368
rect 320234 357312 320956 357368
rect 320173 357310 320956 357312
rect 320173 357307 320239 357310
rect 320950 357308 320956 357310
rect 321020 357308 321026 357372
rect 398925 357370 398991 357373
rect 423121 357372 423187 357373
rect 417182 357370 417188 357372
rect 398925 357368 417188 357370
rect 398925 357312 398930 357368
rect 398986 357312 417188 357368
rect 398925 357310 417188 357312
rect 398925 357307 398991 357310
rect 417182 357308 417188 357310
rect 417252 357308 417258 357372
rect 423070 357370 423076 357372
rect 423030 357310 423076 357370
rect 423140 357368 423187 357372
rect 423182 357312 423187 357368
rect 423070 357308 423076 357310
rect 423140 357308 423187 357312
rect 424542 357308 424548 357372
rect 424612 357370 424618 357372
rect 424961 357370 425027 357373
rect 424612 357368 425027 357370
rect 424612 357312 424966 357368
rect 425022 357312 425027 357368
rect 424612 357310 425027 357312
rect 424612 357308 424618 357310
rect 423121 357307 423187 357308
rect 424961 357307 425027 357310
rect 425421 357372 425487 357373
rect 425421 357368 425468 357372
rect 425532 357370 425538 357372
rect 425421 357312 425426 357368
rect 425421 357308 425468 357312
rect 425532 357310 425578 357370
rect 425532 357308 425538 357310
rect 426566 357308 426572 357372
rect 426636 357370 426642 357372
rect 426893 357370 426959 357373
rect 427629 357372 427695 357373
rect 427629 357370 427676 357372
rect 426636 357368 426959 357370
rect 426636 357312 426898 357368
rect 426954 357312 426959 357368
rect 426636 357310 426959 357312
rect 427584 357368 427676 357370
rect 427584 357312 427634 357368
rect 427584 357310 427676 357312
rect 426636 357308 426642 357310
rect 425421 357307 425487 357308
rect 426893 357307 426959 357310
rect 427629 357308 427676 357310
rect 427740 357308 427746 357372
rect 427813 357370 427879 357373
rect 428549 357372 428615 357373
rect 430021 357372 430087 357373
rect 430573 357372 430639 357373
rect 431953 357372 432019 357373
rect 428222 357370 428228 357372
rect 427813 357368 428228 357370
rect 427813 357312 427818 357368
rect 427874 357312 428228 357368
rect 427813 357310 428228 357312
rect 427629 357307 427695 357308
rect 427813 357307 427879 357310
rect 428222 357308 428228 357310
rect 428292 357308 428298 357372
rect 428549 357368 428596 357372
rect 428660 357370 428666 357372
rect 428549 357312 428554 357368
rect 428549 357308 428596 357312
rect 428660 357310 428706 357370
rect 430021 357368 430068 357372
rect 430132 357370 430138 357372
rect 430573 357370 430620 357372
rect 430021 357312 430026 357368
rect 428660 357308 428666 357310
rect 430021 357308 430068 357312
rect 430132 357310 430178 357370
rect 430528 357368 430620 357370
rect 430528 357312 430578 357368
rect 430528 357310 430620 357312
rect 430132 357308 430138 357310
rect 430573 357308 430620 357310
rect 430684 357308 430690 357372
rect 431902 357308 431908 357372
rect 431972 357370 432019 357372
rect 433333 357370 433399 357373
rect 433558 357370 433564 357372
rect 431972 357368 432064 357370
rect 432014 357312 432064 357368
rect 431972 357310 432064 357312
rect 433333 357368 433564 357370
rect 433333 357312 433338 357368
rect 433394 357312 433564 357368
rect 433333 357310 433564 357312
rect 431972 357308 432019 357310
rect 428549 357307 428615 357308
rect 430021 357307 430087 357308
rect 430573 357307 430639 357308
rect 431953 357307 432019 357308
rect 433333 357307 433399 357310
rect 433558 357308 433564 357310
rect 433628 357308 433634 357372
rect 434713 357370 434779 357373
rect 435950 357370 435956 357372
rect 434713 357368 435956 357370
rect 434713 357312 434718 357368
rect 434774 357312 435956 357368
rect 434713 357310 435956 357312
rect 434713 357307 434779 357310
rect 435950 357308 435956 357310
rect 436020 357308 436026 357372
rect 436829 357370 436895 357373
rect 437054 357370 437060 357372
rect 436829 357368 437060 357370
rect 436829 357312 436834 357368
rect 436890 357312 437060 357368
rect 436829 357310 437060 357312
rect 436829 357307 436895 357310
rect 437054 357308 437060 357310
rect 437124 357308 437130 357372
rect 437473 357370 437539 357373
rect 438526 357370 438532 357372
rect 437473 357368 438532 357370
rect 437473 357312 437478 357368
rect 437534 357312 438532 357368
rect 437473 357310 438532 357312
rect 437473 357307 437539 357310
rect 438526 357308 438532 357310
rect 438596 357308 438602 357372
rect 440233 357370 440299 357373
rect 440918 357370 440924 357372
rect 440233 357368 440924 357370
rect 440233 357312 440238 357368
rect 440294 357312 440924 357368
rect 440233 357310 440924 357312
rect 440233 357307 440299 357310
rect 440918 357308 440924 357310
rect 440988 357308 440994 357372
rect 444281 357370 444347 357373
rect 445845 357372 445911 357373
rect 445845 357370 445892 357372
rect 441570 357368 444347 357370
rect 441570 357312 444286 357368
rect 444342 357312 444347 357368
rect 441570 357310 444347 357312
rect 445800 357368 445892 357370
rect 445800 357312 445850 357368
rect 445800 357310 445892 357312
rect 57094 357172 57100 357236
rect 57164 357234 57170 357236
rect 58617 357234 58683 357237
rect 57164 357232 58683 357234
rect 57164 357176 58622 357232
rect 58678 357176 58683 357232
rect 57164 357174 58683 357176
rect 57164 357172 57170 357174
rect 58617 357171 58683 357174
rect 70710 357172 70716 357236
rect 70780 357234 70786 357236
rect 71589 357234 71655 357237
rect 70780 357232 71655 357234
rect 70780 357176 71594 357232
rect 71650 357176 71655 357232
rect 70780 357174 71655 357176
rect 70780 357172 70786 357174
rect 71589 357171 71655 357174
rect 73286 357172 73292 357236
rect 73356 357234 73362 357236
rect 74073 357234 74139 357237
rect 73356 357232 74139 357234
rect 73356 357176 74078 357232
rect 74134 357176 74139 357232
rect 73356 357174 74139 357176
rect 73356 357172 73362 357174
rect 74073 357171 74139 357174
rect 75862 357172 75868 357236
rect 75932 357234 75938 357236
rect 77017 357234 77083 357237
rect 75932 357232 77083 357234
rect 75932 357176 77022 357232
rect 77078 357176 77083 357232
rect 75932 357174 77083 357176
rect 75932 357172 75938 357174
rect 77017 357171 77083 357174
rect 78254 357172 78260 357236
rect 78324 357234 78330 357236
rect 78489 357234 78555 357237
rect 78324 357232 78555 357234
rect 78324 357176 78494 357232
rect 78550 357176 78555 357232
rect 78324 357174 78555 357176
rect 78324 357172 78330 357174
rect 78489 357171 78555 357174
rect 80646 357172 80652 357236
rect 80716 357234 80722 357236
rect 81249 357234 81315 357237
rect 80716 357232 81315 357234
rect 80716 357176 81254 357232
rect 81310 357176 81315 357232
rect 80716 357174 81315 357176
rect 80716 357172 80722 357174
rect 81249 357171 81315 357174
rect 238017 357234 238083 357237
rect 238334 357234 238340 357236
rect 238017 357232 238340 357234
rect 238017 357176 238022 357232
rect 238078 357176 238340 357232
rect 238017 357174 238340 357176
rect 238017 357171 238083 357174
rect 238334 357172 238340 357174
rect 238404 357234 238410 357236
rect 399385 357234 399451 357237
rect 418102 357234 418108 357236
rect 238404 357232 418108 357234
rect 238404 357176 399390 357232
rect 399446 357176 418108 357232
rect 238404 357174 418108 357176
rect 238404 357172 238410 357174
rect 399385 357171 399451 357174
rect 418102 357172 418108 357174
rect 418172 357172 418178 357236
rect 430665 357234 430731 357237
rect 433425 357236 433491 357237
rect 431166 357234 431172 357236
rect 430665 357232 431172 357234
rect 430665 357176 430670 357232
rect 430726 357176 431172 357232
rect 430665 357174 431172 357176
rect 430665 357171 430731 357174
rect 431166 357172 431172 357174
rect 431236 357172 431242 357236
rect 433374 357234 433380 357236
rect 433334 357174 433380 357234
rect 433444 357232 433491 357236
rect 433486 357176 433491 357232
rect 433374 357172 433380 357174
rect 433444 357172 433491 357176
rect 433425 357171 433491 357172
rect 434621 357236 434687 357237
rect 434621 357232 434668 357236
rect 434732 357234 434738 357236
rect 434621 357176 434626 357232
rect 434621 357172 434668 357176
rect 434732 357174 434778 357234
rect 434732 357172 434738 357174
rect 435766 357172 435772 357236
rect 435836 357234 435842 357236
rect 436001 357234 436067 357237
rect 438393 357236 438459 357237
rect 438342 357234 438348 357236
rect 435836 357232 436067 357234
rect 435836 357176 436006 357232
rect 436062 357176 436067 357232
rect 435836 357174 436067 357176
rect 438302 357174 438348 357234
rect 438412 357232 438459 357236
rect 438454 357176 438459 357232
rect 435836 357172 435842 357174
rect 434621 357171 434687 357172
rect 436001 357171 436067 357174
rect 438342 357172 438348 357174
rect 438412 357172 438459 357176
rect 438894 357172 438900 357236
rect 438964 357234 438970 357236
rect 439446 357234 439452 357236
rect 438964 357174 439452 357234
rect 438964 357172 438970 357174
rect 439446 357172 439452 357174
rect 439516 357234 439522 357236
rect 441570 357234 441630 357310
rect 444281 357307 444347 357310
rect 445845 357308 445892 357310
rect 445956 357308 445962 357372
rect 447225 357370 447291 357373
rect 448278 357370 448284 357372
rect 447225 357368 448284 357370
rect 447225 357312 447230 357368
rect 447286 357312 448284 357368
rect 447225 357310 448284 357312
rect 445845 357307 445911 357308
rect 447225 357307 447291 357310
rect 448278 357308 448284 357310
rect 448348 357308 448354 357372
rect 449893 357370 449959 357373
rect 451038 357370 451044 357372
rect 449893 357368 451044 357370
rect 449893 357312 449898 357368
rect 449954 357312 451044 357368
rect 449893 357310 451044 357312
rect 449893 357307 449959 357310
rect 451038 357308 451044 357310
rect 451108 357308 451114 357372
rect 451457 357370 451523 357373
rect 452142 357370 452148 357372
rect 451457 357368 452148 357370
rect 451457 357312 451462 357368
rect 451518 357312 452148 357368
rect 451457 357310 452148 357312
rect 451457 357307 451523 357310
rect 452142 357308 452148 357310
rect 452212 357308 452218 357372
rect 452653 357370 452719 357373
rect 453614 357370 453620 357372
rect 452653 357368 453620 357370
rect 452653 357312 452658 357368
rect 452714 357312 453620 357368
rect 452653 357310 453620 357312
rect 452653 357307 452719 357310
rect 453614 357308 453620 357310
rect 453684 357308 453690 357372
rect 454677 357370 454743 357373
rect 455822 357370 455828 357372
rect 454677 357368 455828 357370
rect 454677 357312 454682 357368
rect 454738 357312 455828 357368
rect 454677 357310 455828 357312
rect 454677 357307 454743 357310
rect 455822 357308 455828 357310
rect 455892 357308 455898 357372
rect 457529 357370 457595 357373
rect 458398 357370 458404 357372
rect 457529 357368 458404 357370
rect 457529 357312 457534 357368
rect 457590 357312 458404 357368
rect 457529 357310 458404 357312
rect 457529 357307 457595 357310
rect 458398 357308 458404 357310
rect 458468 357308 458474 357372
rect 462313 357370 462379 357373
rect 463550 357370 463556 357372
rect 462313 357368 463556 357370
rect 462313 357312 462318 357368
rect 462374 357312 463556 357368
rect 462313 357310 463556 357312
rect 462313 357307 462379 357310
rect 463550 357308 463556 357310
rect 463620 357308 463626 357372
rect 464337 357370 464403 357373
rect 465942 357370 465948 357372
rect 464337 357368 465948 357370
rect 464337 357312 464342 357368
rect 464398 357312 465948 357368
rect 464337 357310 465948 357312
rect 464337 357307 464403 357310
rect 465942 357308 465948 357310
rect 466012 357308 466018 357372
rect 467833 357370 467899 357373
rect 468150 357370 468156 357372
rect 467833 357368 468156 357370
rect 467833 357312 467838 357368
rect 467894 357312 468156 357368
rect 467833 357310 468156 357312
rect 467833 357307 467899 357310
rect 468150 357308 468156 357310
rect 468220 357308 468226 357372
rect 472617 357370 472683 357373
rect 473302 357370 473308 357372
rect 472617 357368 473308 357370
rect 472617 357312 472622 357368
rect 472678 357312 473308 357368
rect 472617 357310 473308 357312
rect 472617 357307 472683 357310
rect 473302 357308 473308 357310
rect 473372 357308 473378 357372
rect 477493 357370 477559 357373
rect 478454 357370 478460 357372
rect 477493 357368 478460 357370
rect 477493 357312 477498 357368
rect 477554 357312 478460 357368
rect 477493 357310 478460 357312
rect 477493 357307 477559 357310
rect 478454 357308 478460 357310
rect 478524 357308 478530 357372
rect 485773 357370 485839 357373
rect 485998 357370 486004 357372
rect 485773 357368 486004 357370
rect 485773 357312 485778 357368
rect 485834 357312 486004 357368
rect 485773 357310 486004 357312
rect 485773 357307 485839 357310
rect 485998 357308 486004 357310
rect 486068 357308 486074 357372
rect 498193 357370 498259 357373
rect 498510 357370 498516 357372
rect 498193 357368 498516 357370
rect 498193 357312 498198 357368
rect 498254 357312 498516 357368
rect 498193 357310 498516 357312
rect 498193 357307 498259 357310
rect 498510 357308 498516 357310
rect 498580 357308 498586 357372
rect 439516 357174 441630 357234
rect 443085 357234 443151 357237
rect 443494 357234 443500 357236
rect 443085 357232 443500 357234
rect 443085 357176 443090 357232
rect 443146 357176 443500 357232
rect 443085 357174 443500 357176
rect 439516 357172 439522 357174
rect 438393 357171 438459 357172
rect 443085 357171 443151 357174
rect 443494 357172 443500 357174
rect 443564 357172 443570 357236
rect 456793 357234 456859 357237
rect 458030 357234 458036 357236
rect 456793 357232 458036 357234
rect 456793 357176 456798 357232
rect 456854 357176 458036 357232
rect 456793 357174 458036 357176
rect 456793 357171 456859 357174
rect 458030 357172 458036 357174
rect 458100 357172 458106 357236
rect 458173 357234 458239 357237
rect 459134 357234 459140 357236
rect 458173 357232 459140 357234
rect 458173 357176 458178 357232
rect 458234 357176 459140 357232
rect 458173 357174 459140 357176
rect 458173 357171 458239 357174
rect 459134 357172 459140 357174
rect 459204 357172 459210 357236
rect 68318 357036 68324 357100
rect 68388 357098 68394 357100
rect 68921 357098 68987 357101
rect 68388 357096 68987 357098
rect 68388 357040 68926 357096
rect 68982 357040 68987 357096
rect 68388 357038 68987 357040
rect 68388 357036 68394 357038
rect 68921 357035 68987 357038
rect 238753 357098 238819 357101
rect 238886 357098 238892 357100
rect 238753 357096 238892 357098
rect 238753 357040 238758 357096
rect 238814 357040 238892 357096
rect 238753 357038 238892 357040
rect 238753 357035 238819 357038
rect 238886 357036 238892 357038
rect 238956 357098 238962 357100
rect 399569 357098 399635 357101
rect 419574 357098 419580 357100
rect 238956 357096 419580 357098
rect 238956 357040 399574 357096
rect 399630 357040 419580 357096
rect 238956 357038 419580 357040
rect 238956 357036 238962 357038
rect 399569 357035 399635 357038
rect 419574 357036 419580 357038
rect 419644 357036 419650 357100
rect 445661 357098 445727 357101
rect 441570 357096 445727 357098
rect 441570 357040 445666 357096
rect 445722 357040 445727 357096
rect 441570 357038 445727 357040
rect 244590 356900 244596 356964
rect 244660 356962 244666 356964
rect 244917 356962 244983 356965
rect 244660 356960 244983 356962
rect 244660 356904 244922 356960
rect 244978 356904 244983 356960
rect 244660 356902 244983 356904
rect 244660 356900 244666 356902
rect 244917 356899 244983 356902
rect 245101 356962 245167 356965
rect 399661 356962 399727 356965
rect 419942 356962 419948 356964
rect 245101 356960 419948 356962
rect 245101 356904 245106 356960
rect 245162 356904 399666 356960
rect 399722 356904 419948 356960
rect 245101 356902 419948 356904
rect 245101 356899 245167 356902
rect 399661 356899 399727 356902
rect 419942 356900 419948 356902
rect 420012 356900 420018 356964
rect 241830 356826 241836 356828
rect 238710 356766 241836 356826
rect 83590 356628 83596 356692
rect 83660 356690 83666 356692
rect 84101 356690 84167 356693
rect 83660 356688 84167 356690
rect 83660 356632 84106 356688
rect 84162 356632 84167 356688
rect 83660 356630 84167 356632
rect 83660 356628 83666 356630
rect 84101 356627 84167 356630
rect 225229 356690 225295 356693
rect 238710 356690 238770 356766
rect 241830 356764 241836 356766
rect 241900 356826 241906 356828
rect 397177 356826 397243 356829
rect 421782 356826 421788 356828
rect 241900 356824 421788 356826
rect 241900 356768 397182 356824
rect 397238 356768 421788 356824
rect 241900 356766 421788 356768
rect 241900 356764 241906 356766
rect 397177 356763 397243 356766
rect 421782 356764 421788 356766
rect 421852 356764 421858 356828
rect 245561 356692 245627 356693
rect 245510 356690 245516 356692
rect 225229 356688 238770 356690
rect 225229 356632 225234 356688
rect 225290 356632 238770 356688
rect 225229 356630 238770 356632
rect 245470 356630 245516 356690
rect 245580 356688 245627 356692
rect 245622 356632 245627 356688
rect 225229 356627 225295 356630
rect 245510 356628 245516 356630
rect 245580 356628 245627 356632
rect 245561 356627 245627 356628
rect 250069 356692 250135 356693
rect 252277 356692 252343 356693
rect 255773 356692 255839 356693
rect 250069 356688 250116 356692
rect 250180 356690 250186 356692
rect 250069 356632 250074 356688
rect 250069 356628 250116 356632
rect 250180 356630 250226 356690
rect 252277 356688 252324 356692
rect 252388 356690 252394 356692
rect 252277 356632 252282 356688
rect 250180 356628 250186 356630
rect 252277 356628 252324 356632
rect 252388 356630 252434 356690
rect 255773 356688 255820 356692
rect 255884 356690 255890 356692
rect 255773 356632 255778 356688
rect 252388 356628 252394 356630
rect 255773 356628 255820 356632
rect 255884 356630 255930 356690
rect 255884 356628 255890 356630
rect 258390 356628 258396 356692
rect 258460 356690 258466 356692
rect 258809 356690 258875 356693
rect 258460 356688 258875 356690
rect 258460 356632 258814 356688
rect 258870 356632 258875 356688
rect 258460 356630 258875 356632
rect 258460 356628 258466 356630
rect 250069 356627 250135 356628
rect 252277 356627 252343 356628
rect 255773 356627 255839 356628
rect 258809 356627 258875 356630
rect 259494 356628 259500 356692
rect 259564 356690 259570 356692
rect 260189 356690 260255 356693
rect 278078 356690 278084 356692
rect 259564 356688 278084 356690
rect 259564 356632 260194 356688
rect 260250 356632 278084 356688
rect 259564 356630 278084 356632
rect 259564 356628 259570 356630
rect 260189 356627 260255 356630
rect 278078 356628 278084 356630
rect 278148 356690 278154 356692
rect 393957 356690 394023 356693
rect 394509 356690 394575 356693
rect 278148 356688 394575 356690
rect 278148 356632 393962 356688
rect 394018 356632 394514 356688
rect 394570 356632 394575 356688
rect 278148 356630 394575 356632
rect 278148 356628 278154 356630
rect 393957 356627 394023 356630
rect 394509 356627 394575 356630
rect 247125 356554 247191 356557
rect 253381 356556 253447 356557
rect 247534 356554 247540 356556
rect 247125 356552 247540 356554
rect 247125 356496 247130 356552
rect 247186 356496 247540 356552
rect 247125 356494 247540 356496
rect 247125 356491 247191 356494
rect 247534 356492 247540 356494
rect 247604 356492 247610 356556
rect 253381 356552 253428 356556
rect 253492 356554 253498 356556
rect 264973 356554 265039 356557
rect 265934 356554 265940 356556
rect 253381 356496 253386 356552
rect 253381 356492 253428 356496
rect 253492 356494 253538 356554
rect 264973 356552 265940 356554
rect 264973 356496 264978 356552
rect 265034 356496 265940 356552
rect 264973 356494 265940 356496
rect 253492 356492 253498 356494
rect 253381 356491 253447 356492
rect 264973 356491 265039 356494
rect 265934 356492 265940 356494
rect 266004 356492 266010 356556
rect 279182 356554 279188 356556
rect 267690 356494 279188 356554
rect 76046 356356 76052 356420
rect 76116 356418 76122 356420
rect 77201 356418 77267 356421
rect 76116 356416 77267 356418
rect 76116 356360 77206 356416
rect 77262 356360 77267 356416
rect 76116 356358 77267 356360
rect 76116 356356 76122 356358
rect 77201 356355 77267 356358
rect 246614 356356 246620 356420
rect 246684 356418 246690 356420
rect 246849 356418 246915 356421
rect 246684 356416 246915 356418
rect 246684 356360 246854 356416
rect 246910 356360 246915 356416
rect 246684 356358 246915 356360
rect 246684 356356 246690 356358
rect 246849 356355 246915 356358
rect 260097 356418 260163 356421
rect 260598 356418 260604 356420
rect 260097 356416 260604 356418
rect 260097 356360 260102 356416
rect 260158 356360 260604 356416
rect 260097 356358 260604 356360
rect 260097 356355 260163 356358
rect 260598 356356 260604 356358
rect 260668 356418 260674 356420
rect 267690 356418 267750 356494
rect 279182 356492 279188 356494
rect 279252 356554 279258 356556
rect 393865 356554 393931 356557
rect 440734 356554 440740 356556
rect 279252 356552 440740 356554
rect 279252 356496 393870 356552
rect 393926 356496 440740 356552
rect 279252 356494 440740 356496
rect 279252 356492 279258 356494
rect 393865 356491 393931 356494
rect 440734 356492 440740 356494
rect 440804 356554 440810 356556
rect 441570 356554 441630 357038
rect 445661 357035 445727 357038
rect 447133 357098 447199 357101
rect 447542 357098 447548 357100
rect 447133 357096 447548 357098
rect 447133 357040 447138 357096
rect 447194 357040 447548 357096
rect 447133 357038 447548 357040
rect 447133 357035 447199 357038
rect 447542 357036 447548 357038
rect 447612 357036 447618 357100
rect 449985 357098 450051 357101
rect 450854 357098 450860 357100
rect 449985 357096 450860 357098
rect 449985 357040 449990 357096
rect 450046 357040 450860 357096
rect 449985 357038 450860 357040
rect 449985 357035 450051 357038
rect 450854 357036 450860 357038
rect 450924 357036 450930 357100
rect 454033 357098 454099 357101
rect 454350 357098 454356 357100
rect 454033 357096 454356 357098
rect 454033 357040 454038 357096
rect 454094 357040 454356 357096
rect 454033 357038 454356 357040
rect 454033 357035 454099 357038
rect 454350 357036 454356 357038
rect 454420 357036 454426 357100
rect 480529 357098 480595 357101
rect 480662 357098 480668 357100
rect 480529 357096 480668 357098
rect 480529 357040 480534 357096
rect 480590 357040 480668 357096
rect 480529 357038 480668 357040
rect 480529 357035 480595 357038
rect 480662 357036 480668 357038
rect 480732 357036 480738 357100
rect 452745 356962 452811 356965
rect 453246 356962 453252 356964
rect 452745 356960 453252 356962
rect 452745 356904 452750 356960
rect 452806 356904 453252 356960
rect 452745 356902 453252 356904
rect 452745 356899 452811 356902
rect 453246 356900 453252 356902
rect 453316 356900 453322 356964
rect 455413 356962 455479 356965
rect 455638 356962 455644 356964
rect 455413 356960 455644 356962
rect 455413 356904 455418 356960
rect 455474 356904 455644 356960
rect 455413 356902 455644 356904
rect 455413 356899 455479 356902
rect 455638 356900 455644 356902
rect 455708 356900 455714 356964
rect 448513 356828 448579 356829
rect 448462 356764 448468 356828
rect 448532 356826 448579 356828
rect 456793 356826 456859 356829
rect 456926 356826 456932 356828
rect 448532 356824 448624 356826
rect 448574 356768 448624 356824
rect 448532 356766 448624 356768
rect 456793 356824 456932 356826
rect 456793 356768 456798 356824
rect 456854 356768 456932 356824
rect 456793 356766 456932 356768
rect 448532 356764 448579 356766
rect 448513 356763 448579 356764
rect 456793 356763 456859 356766
rect 456926 356764 456932 356766
rect 456996 356764 457002 356828
rect 502333 356826 502399 356829
rect 503294 356826 503300 356828
rect 502333 356824 503300 356826
rect 502333 356768 502338 356824
rect 502394 356768 503300 356824
rect 502333 356766 503300 356768
rect 502333 356763 502399 356766
rect 503294 356764 503300 356766
rect 503364 356764 503370 356828
rect 445753 356690 445819 356693
rect 446254 356690 446260 356692
rect 445753 356688 446260 356690
rect 445753 356632 445758 356688
rect 445814 356632 446260 356688
rect 445753 356630 446260 356632
rect 445753 356627 445819 356630
rect 446254 356628 446260 356630
rect 446324 356628 446330 356692
rect 440804 356494 441630 356554
rect 441705 356554 441771 356557
rect 442022 356554 442028 356556
rect 441705 356552 442028 356554
rect 441705 356496 441710 356552
rect 441766 356496 442028 356552
rect 441705 356494 442028 356496
rect 440804 356492 440810 356494
rect 441705 356491 441771 356494
rect 442022 356492 442028 356494
rect 442092 356492 442098 356556
rect 442993 356554 443059 356557
rect 443862 356554 443868 356556
rect 442993 356552 443868 356554
rect 442993 356496 442998 356552
rect 443054 356496 443868 356552
rect 442993 356494 443868 356496
rect 442993 356491 443059 356494
rect 443862 356492 443868 356494
rect 443932 356492 443938 356556
rect 448513 356554 448579 356557
rect 449750 356554 449756 356556
rect 448513 356552 449756 356554
rect 448513 356496 448518 356552
rect 448574 356496 449756 356552
rect 448513 356494 449756 356496
rect 448513 356491 448579 356494
rect 449750 356492 449756 356494
rect 449820 356492 449826 356556
rect 483013 356554 483079 356557
rect 483422 356554 483428 356556
rect 483013 356552 483428 356554
rect 483013 356496 483018 356552
rect 483074 356496 483428 356552
rect 483013 356494 483428 356496
rect 483013 356491 483079 356494
rect 483422 356492 483428 356494
rect 483492 356492 483498 356556
rect 260668 356358 267750 356418
rect 394509 356418 394575 356421
rect 438894 356418 438900 356420
rect 394509 356416 438900 356418
rect 394509 356360 394514 356416
rect 394570 356360 438900 356416
rect 394509 356358 438900 356360
rect 260668 356356 260674 356358
rect 394509 356355 394575 356358
rect 438894 356356 438900 356358
rect 438964 356356 438970 356420
rect 441981 356418 442047 356421
rect 442758 356418 442764 356420
rect 441981 356416 442764 356418
rect 441981 356360 441986 356416
rect 442042 356360 442764 356416
rect 441981 356358 442764 356360
rect 441981 356355 442047 356358
rect 442758 356356 442764 356358
rect 442828 356356 442834 356420
rect 444373 356418 444439 356421
rect 444782 356418 444788 356420
rect 444373 356416 444788 356418
rect 444373 356360 444378 356416
rect 444434 356360 444788 356416
rect 444373 356358 444788 356360
rect 444373 356355 444439 356358
rect 444782 356356 444788 356358
rect 444852 356356 444858 356420
rect 474733 356418 474799 356421
rect 500953 356420 501019 356421
rect 475878 356418 475884 356420
rect 474733 356416 475884 356418
rect 474733 356360 474738 356416
rect 474794 356360 475884 356416
rect 474733 356358 475884 356360
rect 474733 356355 474799 356358
rect 475878 356356 475884 356358
rect 475948 356356 475954 356420
rect 500902 356356 500908 356420
rect 500972 356418 501019 356420
rect 500972 356416 501064 356418
rect 501014 356360 501064 356416
rect 500972 356358 501064 356360
rect 500972 356356 501019 356358
rect 500953 356355 501019 356356
rect 237005 356282 237071 356285
rect 237230 356282 237236 356284
rect 237005 356280 237236 356282
rect 237005 356224 237010 356280
rect 237066 356224 237236 356280
rect 237005 356222 237236 356224
rect 237005 356219 237071 356222
rect 237230 356220 237236 356222
rect 237300 356282 237306 356284
rect 398925 356282 398991 356285
rect 237300 356280 398991 356282
rect 237300 356224 398930 356280
rect 398986 356224 398991 356280
rect 237300 356222 398991 356224
rect 237300 356220 237306 356222
rect 398925 356219 398991 356222
rect 470777 356282 470843 356285
rect 470910 356282 470916 356284
rect 470777 356280 470916 356282
rect 470777 356224 470782 356280
rect 470838 356224 470916 356280
rect 470777 356222 470916 356224
rect 470777 356219 470843 356222
rect 470910 356220 470916 356222
rect 470980 356220 470986 356284
rect 489678 356220 489684 356284
rect 489748 356282 489754 356284
rect 489913 356282 489979 356285
rect 489748 356280 489979 356282
rect 489748 356224 489918 356280
rect 489974 356224 489979 356280
rect 489748 356222 489979 356224
rect 489748 356220 489754 356222
rect 489913 356219 489979 356222
rect 495433 356282 495499 356285
rect 495566 356282 495572 356284
rect 495433 356280 495572 356282
rect 495433 356224 495438 356280
rect 495494 356224 495572 356280
rect 495433 356222 495572 356224
rect 495433 356219 495499 356222
rect 495566 356220 495572 356222
rect 495636 356220 495642 356284
rect 64638 356084 64644 356148
rect 64708 356146 64714 356148
rect 66161 356146 66227 356149
rect 64708 356144 66227 356146
rect 64708 356088 66166 356144
rect 66222 356088 66227 356144
rect 64708 356086 66227 356088
rect 64708 356084 64714 356086
rect 66161 356083 66227 356086
rect 67582 356084 67588 356148
rect 67652 356146 67658 356148
rect 68921 356146 68987 356149
rect 67652 356144 68987 356146
rect 67652 356088 68926 356144
rect 68982 356088 68987 356144
rect 67652 356086 68987 356088
rect 67652 356084 67658 356086
rect 68921 356083 68987 356086
rect 103278 356084 103284 356148
rect 103348 356146 103354 356148
rect 104801 356146 104867 356149
rect 103348 356144 104867 356146
rect 103348 356088 104806 356144
rect 104862 356088 104867 356144
rect 103348 356086 104867 356088
rect 103348 356084 103354 356086
rect 104801 356083 104867 356086
rect 240910 356084 240916 356148
rect 240980 356084 240986 356148
rect 245101 356146 245167 356149
rect 241470 356144 245167 356146
rect 241470 356088 245106 356144
rect 245162 356088 245167 356144
rect 241470 356086 245167 356088
rect 213269 356010 213335 356013
rect 240225 356010 240291 356013
rect 240918 356010 240978 356084
rect 241470 356010 241530 356086
rect 245101 356083 245167 356086
rect 273345 356146 273411 356149
rect 273478 356146 273484 356148
rect 273345 356144 273484 356146
rect 273345 356088 273350 356144
rect 273406 356088 273484 356144
rect 273345 356086 273484 356088
rect 273345 356083 273411 356086
rect 273478 356084 273484 356086
rect 273548 356084 273554 356148
rect 277393 356146 277459 356149
rect 278446 356146 278452 356148
rect 277393 356144 278452 356146
rect 277393 356088 277398 356144
rect 277454 356088 278452 356144
rect 277393 356086 278452 356088
rect 277393 356083 277459 356086
rect 278446 356084 278452 356086
rect 278516 356084 278522 356148
rect 280153 356146 280219 356149
rect 280838 356146 280844 356148
rect 280153 356144 280844 356146
rect 280153 356088 280158 356144
rect 280214 356088 280844 356144
rect 280153 356086 280844 356088
rect 280153 356083 280219 356086
rect 280838 356084 280844 356086
rect 280908 356084 280914 356148
rect 322933 356146 322999 356149
rect 460933 356148 460999 356149
rect 323342 356146 323348 356148
rect 322933 356144 323348 356146
rect 322933 356088 322938 356144
rect 322994 356088 323348 356144
rect 322933 356086 323348 356088
rect 322933 356083 322999 356086
rect 323342 356084 323348 356086
rect 323412 356084 323418 356148
rect 460933 356144 460980 356148
rect 461044 356146 461050 356148
rect 492673 356146 492739 356149
rect 493358 356146 493364 356148
rect 460933 356088 460938 356144
rect 460933 356084 460980 356088
rect 461044 356086 461090 356146
rect 492673 356144 493364 356146
rect 492673 356088 492678 356144
rect 492734 356088 493364 356144
rect 492673 356086 493364 356088
rect 461044 356084 461050 356086
rect 460933 356083 460999 356084
rect 492673 356083 492739 356086
rect 493358 356084 493364 356086
rect 493428 356084 493434 356148
rect 505093 356146 505159 356149
rect 505502 356146 505508 356148
rect 505093 356144 505508 356146
rect 505093 356088 505098 356144
rect 505154 356088 505508 356144
rect 505093 356086 505508 356088
rect 505093 356083 505159 356086
rect 505502 356084 505508 356086
rect 505572 356084 505578 356148
rect 213269 356008 241530 356010
rect 213269 355952 213274 356008
rect 213330 355952 240230 356008
rect 240286 355952 241530 356008
rect 213269 355950 241530 355952
rect 213269 355947 213335 355950
rect 240225 355947 240291 355950
rect 213637 355874 213703 355877
rect 236269 355874 236335 355877
rect 213637 355872 236335 355874
rect 213637 355816 213642 355872
rect 213698 355816 236274 355872
rect 236330 355816 236335 355872
rect 213637 355814 236335 355816
rect 213637 355811 213703 355814
rect 236269 355811 236335 355814
rect 213729 355738 213795 355741
rect 240317 355738 240383 355741
rect 213729 355736 240383 355738
rect 213729 355680 213734 355736
rect 213790 355680 240322 355736
rect 240378 355680 240383 355736
rect 213729 355678 240383 355680
rect 213729 355675 213795 355678
rect 240317 355675 240383 355678
rect 213821 355602 213887 355605
rect 243997 355602 244063 355605
rect 213821 355600 244063 355602
rect 213821 355544 213826 355600
rect 213882 355544 244002 355600
rect 244058 355544 244063 355600
rect 213821 355542 244063 355544
rect 213821 355539 213887 355542
rect 243997 355539 244063 355542
rect 215150 355404 215156 355468
rect 215220 355466 215226 355468
rect 247309 355466 247375 355469
rect 215220 355464 247375 355466
rect 215220 355408 247314 355464
rect 247370 355408 247375 355464
rect 215220 355406 247375 355408
rect 215220 355404 215226 355406
rect 247309 355403 247375 355406
rect 144637 355330 144703 355333
rect 215886 355330 215892 355332
rect 144637 355328 215892 355330
rect 144637 355272 144642 355328
rect 144698 355272 215892 355328
rect 144637 355270 215892 355272
rect 144637 355267 144703 355270
rect 215886 355268 215892 355270
rect 215956 355268 215962 355332
rect 274173 354514 274239 354517
rect 398465 354514 398531 354517
rect 274173 354512 398531 354514
rect 274173 354456 274178 354512
rect 274234 354456 398470 354512
rect 398526 354456 398531 354512
rect 274173 354454 398531 354456
rect 274173 354451 274239 354454
rect 398465 354451 398531 354454
rect 267917 354378 267983 354381
rect 397913 354378 397979 354381
rect 267917 354376 397979 354378
rect 267917 354320 267922 354376
rect 267978 354320 397918 354376
rect 397974 354320 397979 354376
rect 267917 354318 397979 354320
rect 267917 354315 267983 354318
rect 397913 354315 397979 354318
rect 257981 354242 258047 354245
rect 398281 354242 398347 354245
rect 257981 354240 398347 354242
rect 257981 354184 257986 354240
rect 258042 354184 398286 354240
rect 398342 354184 398347 354240
rect 257981 354182 398347 354184
rect 257981 354179 258047 354182
rect 398281 354179 398347 354182
rect 251357 354106 251423 354109
rect 398097 354106 398163 354109
rect 251357 354104 398163 354106
rect 251357 354048 251362 354104
rect 251418 354048 398102 354104
rect 398158 354048 398163 354104
rect 251357 354046 398163 354048
rect 251357 354043 251423 354046
rect 398097 354043 398163 354046
rect 138749 353970 138815 353973
rect 580349 353970 580415 353973
rect 138749 353968 580415 353970
rect 138749 353912 138754 353968
rect 138810 353912 580354 353968
rect 580410 353912 580415 353968
rect 138749 353910 580415 353912
rect 138749 353907 138815 353910
rect 580349 353907 580415 353910
rect 142797 352610 142863 352613
rect 397494 352610 397500 352612
rect 142797 352608 397500 352610
rect 142797 352552 142802 352608
rect 142858 352552 397500 352608
rect 142797 352550 397500 352552
rect 142797 352547 142863 352550
rect 397494 352548 397500 352550
rect 397564 352548 397570 352612
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 255037 351386 255103 351389
rect 392669 351386 392735 351389
rect 255037 351384 392735 351386
rect 255037 351328 255042 351384
rect 255098 351328 392674 351384
rect 392730 351328 392735 351384
rect 255037 351326 392735 351328
rect 255037 351323 255103 351326
rect 392669 351323 392735 351326
rect 237005 351250 237071 351253
rect 399518 351250 399524 351252
rect 237005 351248 399524 351250
rect 237005 351192 237010 351248
rect 237066 351192 399524 351248
rect 237005 351190 399524 351192
rect 237005 351187 237071 351190
rect 399518 351188 399524 351190
rect 399588 351188 399594 351252
rect 141325 351114 141391 351117
rect 395286 351114 395292 351116
rect 141325 351112 395292 351114
rect 141325 351056 141330 351112
rect 141386 351056 395292 351112
rect 141325 351054 395292 351056
rect 141325 351051 141391 351054
rect 395286 351052 395292 351054
rect 395356 351052 395362 351116
rect 140589 349754 140655 349757
rect 398598 349754 398604 349756
rect 140589 349752 398604 349754
rect 140589 349696 140594 349752
rect 140650 349696 398604 349752
rect 140589 349694 398604 349696
rect 140589 349691 140655 349694
rect 398598 349692 398604 349694
rect 398668 349692 398674 349756
rect 237373 348394 237439 348397
rect 399334 348394 399340 348396
rect 237373 348392 399340 348394
rect 237373 348336 237378 348392
rect 237434 348336 399340 348392
rect 237373 348334 399340 348336
rect 237373 348331 237439 348334
rect 399334 348332 399340 348334
rect 399404 348332 399410 348396
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 145005 342954 145071 342957
rect 211654 342954 211660 342956
rect 145005 342952 211660 342954
rect 145005 342896 145010 342952
rect 145066 342896 211660 342952
rect 145005 342894 211660 342896
rect 145005 342891 145071 342894
rect 211654 342892 211660 342894
rect 211724 342892 211730 342956
rect 217358 342892 217364 342956
rect 217428 342954 217434 342956
rect 316677 342954 316743 342957
rect 217428 342952 316743 342954
rect 217428 342896 316682 342952
rect 316738 342896 316743 342952
rect 217428 342894 316743 342896
rect 217428 342892 217434 342894
rect 316677 342891 316743 342894
rect 583520 338452 584960 338692
rect 143901 337378 143967 337381
rect 213126 337378 213132 337380
rect 143901 337376 213132 337378
rect 143901 337320 143906 337376
rect 143962 337320 213132 337376
rect 143901 337318 213132 337320
rect 143901 337315 143967 337318
rect 213126 337316 213132 337318
rect 213196 337316 213202 337380
rect -960 332196 480 332436
rect 145741 327722 145807 327725
rect 214414 327722 214420 327724
rect 145741 327720 214420 327722
rect 145741 327664 145746 327720
rect 145802 327664 214420 327720
rect 145741 327662 214420 327664
rect 145741 327659 145807 327662
rect 214414 327660 214420 327662
rect 214484 327660 214490 327724
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 38694 324940 38700 325004
rect 38764 325002 38770 325004
rect 234429 325002 234495 325005
rect 38764 325000 234495 325002
rect 38764 324944 234434 325000
rect 234490 324944 234495 325000
rect 38764 324942 234495 324944
rect 38764 324940 38770 324942
rect 234429 324939 234495 324942
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 220077 311130 220143 311133
rect 398782 311130 398788 311132
rect 220077 311128 398788 311130
rect 220077 311072 220082 311128
rect 220138 311072 398788 311128
rect 220077 311070 398788 311072
rect 220077 311067 220143 311070
rect 398782 311068 398788 311070
rect 398852 311068 398858 311132
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 38878 304132 38884 304196
rect 38948 304194 38954 304196
rect 238477 304194 238543 304197
rect 38948 304192 238543 304194
rect 38948 304136 238482 304192
rect 238538 304136 238543 304192
rect 38948 304134 238543 304136
rect 38948 304132 38954 304134
rect 238477 304131 238543 304134
rect 229277 298754 229343 298757
rect 357014 298754 357020 298756
rect 229277 298752 357020 298754
rect 229277 298696 229282 298752
rect 229338 298696 357020 298752
rect 229277 298694 357020 298696
rect 229277 298691 229343 298694
rect 357014 298692 357020 298694
rect 357084 298692 357090 298756
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 233325 297394 233391 297397
rect 356646 297394 356652 297396
rect 233325 297392 356652 297394
rect 233325 297336 233330 297392
rect 233386 297336 356652 297392
rect 233325 297334 356652 297336
rect 233325 297331 233391 297334
rect 356646 297332 356652 297334
rect 356716 297332 356722 297396
rect 208669 294538 208735 294541
rect 357934 294538 357940 294540
rect 208669 294536 357940 294538
rect 208669 294480 208674 294536
rect 208730 294480 357940 294536
rect 208669 294478 357940 294480
rect 208669 294475 208735 294478
rect 357934 294476 357940 294478
rect 358004 294476 358010 294540
rect 206318 293524 206324 293588
rect 206388 293586 206394 293588
rect 249517 293586 249583 293589
rect 206388 293584 249583 293586
rect 206388 293528 249522 293584
rect 249578 293528 249583 293584
rect 206388 293526 249583 293528
rect 206388 293524 206394 293526
rect 249517 293523 249583 293526
rect 206134 293388 206140 293452
rect 206204 293450 206210 293452
rect 292941 293450 293007 293453
rect 206204 293448 293007 293450
rect 206204 293392 292946 293448
rect 293002 293392 293007 293448
rect 206204 293390 293007 293392
rect 206204 293388 206210 293390
rect 292941 293387 293007 293390
rect -960 293178 480 293268
rect 203374 293252 203380 293316
rect 203444 293314 203450 293316
rect 313549 293314 313615 293317
rect 203444 293312 313615 293314
rect 203444 293256 313554 293312
rect 313610 293256 313615 293312
rect 203444 293254 313615 293256
rect 203444 293252 203450 293254
rect 313549 293251 313615 293254
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 213085 293178 213151 293181
rect 359406 293178 359412 293180
rect 213085 293176 359412 293178
rect 213085 293120 213090 293176
rect 213146 293120 359412 293176
rect 213085 293118 359412 293120
rect 213085 293115 213151 293118
rect 359406 293116 359412 293118
rect 359476 293116 359482 293180
rect 203609 291002 203675 291005
rect 227069 291002 227135 291005
rect 203609 291000 227135 291002
rect 203609 290944 203614 291000
rect 203670 290944 227074 291000
rect 227130 290944 227135 291000
rect 203609 290942 227135 290944
rect 203609 290939 203675 290942
rect 227069 290939 227135 290942
rect 177481 290866 177547 290869
rect 252829 290866 252895 290869
rect 177481 290864 252895 290866
rect 177481 290808 177486 290864
rect 177542 290808 252834 290864
rect 252890 290808 252895 290864
rect 177481 290806 252895 290808
rect 177481 290803 177547 290806
rect 252829 290803 252895 290806
rect 177665 290730 177731 290733
rect 256141 290730 256207 290733
rect 177665 290728 256207 290730
rect 177665 290672 177670 290728
rect 177726 290672 256146 290728
rect 256202 290672 256207 290728
rect 177665 290670 256207 290672
rect 177665 290667 177731 290670
rect 256141 290667 256207 290670
rect 140957 290594 141023 290597
rect 542353 290594 542419 290597
rect 140957 290592 542419 290594
rect 140957 290536 140962 290592
rect 141018 290536 542358 290592
rect 542414 290536 542419 290592
rect 140957 290534 542419 290536
rect 140957 290531 141023 290534
rect 542353 290531 542419 290534
rect 133965 290458 134031 290461
rect 548517 290458 548583 290461
rect 133965 290456 548583 290458
rect 133965 290400 133970 290456
rect 134026 290400 548522 290456
rect 548578 290400 548583 290456
rect 133965 290398 548583 290400
rect 133965 290395 134031 290398
rect 548517 290395 548583 290398
rect 219934 289036 219940 289100
rect 220004 289098 220010 289100
rect 262765 289098 262831 289101
rect 220004 289096 262831 289098
rect 220004 289040 262770 289096
rect 262826 289040 262831 289096
rect 220004 289038 262831 289040
rect 220004 289036 220010 289038
rect 262765 289035 262831 289038
rect 214598 287812 214604 287876
rect 214668 287874 214674 287876
rect 269021 287874 269087 287877
rect 214668 287872 269087 287874
rect 214668 287816 269026 287872
rect 269082 287816 269087 287872
rect 214668 287814 269087 287816
rect 214668 287812 214674 287814
rect 269021 287811 269087 287814
rect 214782 287676 214788 287740
rect 214852 287738 214858 287740
rect 271965 287738 272031 287741
rect 214852 287736 272031 287738
rect 214852 287680 271970 287736
rect 272026 287680 272031 287736
rect 214852 287678 272031 287680
rect 214852 287676 214858 287678
rect 271965 287675 272031 287678
rect 189901 287466 189967 287469
rect 319621 287466 319687 287469
rect 189901 287464 319687 287466
rect 189901 287408 189906 287464
rect 189962 287408 319626 287464
rect 319682 287408 319687 287464
rect 189901 287406 319687 287408
rect 189901 287403 189967 287406
rect 319621 287403 319687 287406
rect 181805 287330 181871 287333
rect 320817 287330 320883 287333
rect 181805 287328 320883 287330
rect 181805 287272 181810 287328
rect 181866 287272 320822 287328
rect 320878 287272 320883 287328
rect 181805 287270 320883 287272
rect 181805 287267 181871 287270
rect 320817 287267 320883 287270
rect 187693 287194 187759 287197
rect 517513 287194 517579 287197
rect 187693 287192 517579 287194
rect 187693 287136 187698 287192
rect 187754 287136 517518 287192
rect 517574 287136 517579 287192
rect 187693 287134 517579 287136
rect 187693 287131 187759 287134
rect 517513 287131 517579 287134
rect 214741 285426 214807 285429
rect 255589 285426 255655 285429
rect 214741 285424 255655 285426
rect 214741 285368 214746 285424
rect 214802 285368 255594 285424
rect 255650 285368 255655 285424
rect 214741 285366 255655 285368
rect 214741 285363 214807 285366
rect 255589 285363 255655 285366
rect 214281 285290 214347 285293
rect 258901 285290 258967 285293
rect 214281 285288 258967 285290
rect 214281 285232 214286 285288
rect 214342 285232 258906 285288
rect 258962 285232 258967 285288
rect 583520 285276 584960 285516
rect 214281 285230 258967 285232
rect 214281 285227 214347 285230
rect 258901 285227 258967 285230
rect 214465 285154 214531 285157
rect 262213 285154 262279 285157
rect 214465 285152 262279 285154
rect 214465 285096 214470 285152
rect 214526 285096 262218 285152
rect 262274 285096 262279 285152
rect 214465 285094 262279 285096
rect 214465 285091 214531 285094
rect 262213 285091 262279 285094
rect 215017 285018 215083 285021
rect 265525 285018 265591 285021
rect 215017 285016 265591 285018
rect 215017 284960 215022 285016
rect 215078 284960 265530 285016
rect 265586 284960 265591 285016
rect 215017 284958 265591 284960
rect 215017 284955 215083 284958
rect 265525 284955 265591 284958
rect 136449 284882 136515 284885
rect 544377 284882 544443 284885
rect 136449 284880 544443 284882
rect 136449 284824 136454 284880
rect 136510 284824 544382 284880
rect 544438 284824 544443 284880
rect 136449 284822 544443 284824
rect 136449 284819 136515 284822
rect 544377 284819 544443 284822
rect 178125 282842 178191 282845
rect 161430 282840 178191 282842
rect 161430 282784 178130 282840
rect 178186 282784 178191 282840
rect 161430 282782 178191 282784
rect 148593 282162 148659 282165
rect 161430 282162 161490 282782
rect 178125 282779 178191 282782
rect 208710 282780 208716 282844
rect 208780 282842 208786 282844
rect 209221 282842 209287 282845
rect 208780 282840 209287 282842
rect 208780 282784 209226 282840
rect 209282 282784 209287 282840
rect 208780 282782 209287 282784
rect 208780 282780 208786 282782
rect 209221 282779 209287 282782
rect 210693 282842 210759 282845
rect 210918 282842 210924 282844
rect 210693 282840 210924 282842
rect 210693 282784 210698 282840
rect 210754 282784 210924 282840
rect 210693 282782 210924 282784
rect 210693 282779 210759 282782
rect 210918 282780 210924 282782
rect 210988 282780 210994 282844
rect 211521 282842 211587 282845
rect 212206 282842 212212 282844
rect 211521 282840 212212 282842
rect 211521 282784 211526 282840
rect 211582 282784 212212 282840
rect 211521 282782 212212 282784
rect 211521 282779 211587 282782
rect 212206 282780 212212 282782
rect 212276 282780 212282 282844
rect 215845 282842 215911 282845
rect 216070 282842 216076 282844
rect 215845 282840 216076 282842
rect 215845 282784 215850 282840
rect 215906 282784 216076 282840
rect 215845 282782 216076 282784
rect 215845 282779 215911 282782
rect 216070 282780 216076 282782
rect 216140 282780 216146 282844
rect 216213 282842 216279 282845
rect 216438 282842 216444 282844
rect 216213 282840 216444 282842
rect 216213 282784 216218 282840
rect 216274 282784 216444 282840
rect 216213 282782 216444 282784
rect 216213 282779 216279 282782
rect 216438 282780 216444 282782
rect 216508 282780 216514 282844
rect 216622 282780 216628 282844
rect 216692 282842 216698 282844
rect 217685 282842 217751 282845
rect 216692 282840 217751 282842
rect 216692 282784 217690 282840
rect 217746 282784 217751 282840
rect 216692 282782 217751 282784
rect 216692 282780 216698 282782
rect 217685 282779 217751 282782
rect 218421 282842 218487 282845
rect 218646 282842 218652 282844
rect 218421 282840 218652 282842
rect 218421 282784 218426 282840
rect 218482 282784 218652 282840
rect 218421 282782 218652 282784
rect 218421 282779 218487 282782
rect 218646 282780 218652 282782
rect 218716 282780 218722 282844
rect 219750 282780 219756 282844
rect 219820 282842 219826 282844
rect 220261 282842 220327 282845
rect 219820 282840 220327 282842
rect 219820 282784 220266 282840
rect 220322 282784 220327 282840
rect 219820 282782 220327 282784
rect 219820 282780 219826 282782
rect 220261 282779 220327 282782
rect 211613 282706 211679 282709
rect 212390 282706 212396 282708
rect 211613 282704 212396 282706
rect 211613 282648 211618 282704
rect 211674 282648 212396 282704
rect 211613 282646 212396 282648
rect 211613 282643 211679 282646
rect 212390 282644 212396 282646
rect 212460 282644 212466 282708
rect 212574 282644 212580 282708
rect 212644 282706 212650 282708
rect 213637 282706 213703 282709
rect 212644 282704 213703 282706
rect 212644 282648 213642 282704
rect 213698 282648 213703 282704
rect 212644 282646 213703 282648
rect 212644 282644 212650 282646
rect 213637 282643 213703 282646
rect 217542 282508 217548 282572
rect 217612 282570 217618 282572
rect 248965 282570 249031 282573
rect 217612 282568 249031 282570
rect 217612 282512 248970 282568
rect 249026 282512 249031 282568
rect 217612 282510 249031 282512
rect 217612 282508 217618 282510
rect 248965 282507 249031 282510
rect 315757 282298 315823 282301
rect 358118 282298 358124 282300
rect 315757 282296 358124 282298
rect 315757 282240 315762 282296
rect 315818 282240 358124 282296
rect 315757 282238 358124 282240
rect 315757 282235 315823 282238
rect 358118 282236 358124 282238
rect 358188 282236 358194 282300
rect 148593 282160 161490 282162
rect 148593 282104 148598 282160
rect 148654 282104 161490 282160
rect 148593 282102 161490 282104
rect 183461 282162 183527 282165
rect 319805 282162 319871 282165
rect 183461 282160 319871 282162
rect 183461 282104 183466 282160
rect 183522 282104 319810 282160
rect 319866 282104 319871 282160
rect 183461 282102 319871 282104
rect 148593 282099 148659 282102
rect 183461 282099 183527 282102
rect 319805 282099 319871 282102
rect 188981 282026 189047 282029
rect 456057 282026 456123 282029
rect 188981 282024 456123 282026
rect 188981 281968 188986 282024
rect 189042 281968 456062 282024
rect 456118 281968 456123 282024
rect 188981 281966 456123 281968
rect 188981 281963 189047 281966
rect 456057 281963 456123 281966
rect 126881 281890 126947 281893
rect 175181 281890 175247 281893
rect 126881 281888 175247 281890
rect 126881 281832 126886 281888
rect 126942 281832 175186 281888
rect 175242 281832 175247 281888
rect 126881 281830 175247 281832
rect 126881 281827 126947 281830
rect 175181 281827 175247 281830
rect 191281 281890 191347 281893
rect 469857 281890 469923 281893
rect 191281 281888 469923 281890
rect 191281 281832 191286 281888
rect 191342 281832 469862 281888
rect 469918 281832 469923 281888
rect 191281 281830 469923 281832
rect 191281 281827 191347 281830
rect 469857 281827 469923 281830
rect 125501 281754 125567 281757
rect 175917 281754 175983 281757
rect 125501 281752 175983 281754
rect 125501 281696 125506 281752
rect 125562 281696 175922 281752
rect 175978 281696 175983 281752
rect 125501 281694 175983 281696
rect 125501 281691 125567 281694
rect 175917 281691 175983 281694
rect 178769 281754 178835 281757
rect 491937 281754 492003 281757
rect 178769 281752 492003 281754
rect 178769 281696 178774 281752
rect 178830 281696 491942 281752
rect 491998 281696 492003 281752
rect 178769 281694 492003 281696
rect 178769 281691 178835 281694
rect 491937 281691 492003 281694
rect 128721 281618 128787 281621
rect 185577 281618 185643 281621
rect 128721 281616 185643 281618
rect 128721 281560 128726 281616
rect 128782 281560 185582 281616
rect 185638 281560 185643 281616
rect 128721 281558 185643 281560
rect 128721 281555 128787 281558
rect 185577 281555 185643 281558
rect 186221 281618 186287 281621
rect 514753 281618 514819 281621
rect 186221 281616 514819 281618
rect 186221 281560 186226 281616
rect 186282 281560 514758 281616
rect 514814 281560 514819 281616
rect 186221 281558 514819 281560
rect 186221 281555 186287 281558
rect 514753 281555 514819 281558
rect 175917 280938 175983 280941
rect 580257 280938 580323 280941
rect 175917 280936 580323 280938
rect 175917 280880 175922 280936
rect 175978 280880 580262 280936
rect 580318 280880 580323 280936
rect 175917 280878 580323 280880
rect 175917 280875 175983 280878
rect 580257 280875 580323 280878
rect 175181 280802 175247 280805
rect 580441 280802 580507 280805
rect 175181 280800 580507 280802
rect 175181 280744 175186 280800
rect 175242 280744 580446 280800
rect 580502 280744 580507 280800
rect 175181 280742 580507 280744
rect 175181 280739 175247 280742
rect 580441 280739 580507 280742
rect 127755 280258 127821 280261
rect 540329 280258 540395 280261
rect 127755 280256 540395 280258
rect -960 279972 480 280212
rect 127755 280200 127760 280256
rect 127816 280200 540334 280256
rect 540390 280200 540395 280256
rect 127755 280198 540395 280200
rect 127755 280195 127821 280198
rect 540329 280195 540395 280198
rect 123702 279516 123708 279580
rect 123772 279578 123778 279580
rect 123845 279578 123911 279581
rect 123772 279576 123911 279578
rect 123772 279520 123850 279576
rect 123906 279520 123911 279576
rect 123772 279518 123911 279520
rect 123772 279516 123778 279518
rect 123845 279515 123911 279518
rect 123707 279306 123773 279309
rect 123886 279306 123892 279308
rect 123707 279304 123892 279306
rect 123707 279248 123712 279304
rect 123768 279248 123892 279304
rect 123707 279246 123892 279248
rect 123707 279243 123773 279246
rect 123886 279244 123892 279246
rect 123956 279244 123962 279308
rect 583520 272234 584960 272324
rect 567150 272174 584960 272234
rect 318241 271962 318307 271965
rect 567150 271962 567210 272174
rect 583520 272084 584960 272174
rect 318241 271960 567210 271962
rect 318241 271904 318246 271960
rect 318302 271904 567210 271960
rect 318241 271902 567210 271904
rect 318241 271899 318307 271902
rect -960 267202 480 267292
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2957 254146 3023 254149
rect -960 254144 3023 254146
rect -960 254088 2962 254144
rect 3018 254088 3023 254144
rect -960 254086 3023 254088
rect -960 253996 480 254086
rect 2957 254083 3023 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 318149 233882 318215 233885
rect 498929 233882 498995 233885
rect 318149 233880 498995 233882
rect 318149 233824 318154 233880
rect 318210 233824 498934 233880
rect 498990 233824 498995 233880
rect 318149 233822 498995 233824
rect 318149 233819 318215 233822
rect 498929 233819 498995 233822
rect 318057 232522 318123 232525
rect 513281 232522 513347 232525
rect 318057 232520 513347 232522
rect 318057 232464 318062 232520
rect 318118 232464 513286 232520
rect 513342 232464 513347 232520
rect 318057 232462 513347 232464
rect 318057 232459 318123 232462
rect 513281 232459 513347 232462
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 318057 230618 318123 230621
rect 534809 230618 534875 230621
rect 318057 230616 534875 230618
rect 318057 230560 318062 230616
rect 318118 230560 534814 230616
rect 534870 230560 534875 230616
rect 318057 230558 534875 230560
rect 318057 230555 318123 230558
rect 534809 230555 534875 230558
rect 532417 229258 532483 229261
rect 528510 229256 532483 229258
rect 528510 229200 532422 229256
rect 532478 229200 532483 229256
rect 528510 229198 532483 229200
rect 318149 229122 318215 229125
rect 528510 229122 528570 229198
rect 532417 229195 532483 229198
rect 318149 229120 528570 229122
rect 318149 229064 318154 229120
rect 318210 229064 528570 229120
rect 318149 229062 528570 229064
rect 318149 229059 318215 229062
rect -960 227884 480 228124
rect 580717 219058 580783 219061
rect 583520 219058 584960 219148
rect 580717 219056 584960 219058
rect 580717 219000 580722 219056
rect 580778 219000 584960 219056
rect 580717 218998 584960 219000
rect 580717 218995 580783 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3049 214978 3115 214981
rect -960 214976 3115 214978
rect -960 214920 3054 214976
rect 3110 214920 3115 214976
rect -960 214918 3115 214920
rect -960 214828 480 214918
rect 3049 214915 3115 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3785 201922 3851 201925
rect -960 201920 3851 201922
rect -960 201864 3790 201920
rect 3846 201864 3851 201920
rect -960 201862 3851 201864
rect -960 201772 480 201862
rect 3785 201859 3851 201862
rect 580625 192538 580691 192541
rect 583520 192538 584960 192628
rect 580625 192536 584960 192538
rect 580625 192480 580630 192536
rect 580686 192480 584960 192536
rect 580625 192478 584960 192480
rect 580625 192475 580691 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 580533 179210 580599 179213
rect 583520 179210 584960 179300
rect 580533 179208 584960 179210
rect 580533 179152 580538 179208
rect 580594 179152 584960 179208
rect 580533 179150 584960 179152
rect 580533 179147 580599 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3049 162890 3115 162893
rect -960 162888 3115 162890
rect -960 162832 3054 162888
rect 3110 162832 3115 162888
rect -960 162830 3115 162832
rect -960 162740 480 162830
rect 3049 162827 3115 162830
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 580349 152627 580415 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 579797 139362 579863 139365
rect 583520 139362 584960 139452
rect 579797 139360 584960 139362
rect 579797 139304 579802 139360
rect 579858 139304 584960 139360
rect 579797 139302 584960 139304
rect 579797 139299 579863 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579613 112842 579679 112845
rect 583520 112842 584960 112932
rect 579613 112840 584960 112842
rect 579613 112784 579618 112840
rect 579674 112784 584960 112840
rect 579613 112782 584960 112784
rect 579613 112779 579679 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 580441 99514 580507 99517
rect 583520 99514 584960 99604
rect 580441 99512 584960 99514
rect 580441 99456 580446 99512
rect 580502 99456 584960 99512
rect 580441 99454 584960 99456
rect 580441 99451 580507 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3325 97610 3391 97613
rect -960 97608 3391 97610
rect -960 97552 3330 97608
rect 3386 97552 3391 97608
rect -960 97550 3391 97552
rect -960 97460 480 97550
rect 3325 97547 3391 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3693 84690 3759 84693
rect -960 84688 3759 84690
rect -960 84632 3698 84688
rect 3754 84632 3759 84688
rect -960 84630 3759 84632
rect -960 84540 480 84630
rect 3693 84627 3759 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3601 71634 3667 71637
rect -960 71632 3667 71634
rect -960 71576 3606 71632
rect 3662 71576 3667 71632
rect -960 71574 3667 71576
rect -960 71484 480 71574
rect 3601 71571 3667 71574
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 123702 31724 123708 31788
rect 123772 31786 123778 31788
rect 583526 31786 583586 32950
rect 123772 31726 583586 31786
rect 123772 31724 123778 31726
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 123886 7516 123892 7580
rect 123956 7578 123962 7580
rect 579981 7578 580047 7581
rect 123956 7576 580047 7578
rect 123956 7520 579986 7576
rect 580042 7520 580047 7576
rect 123956 7518 580047 7520
rect 123956 7516 123962 7518
rect 579981 7515 580047 7518
rect 579981 6626 580047 6629
rect 583520 6626 584960 6716
rect 579981 6624 584960 6626
rect -960 6490 480 6580
rect 579981 6568 579986 6624
rect 580042 6568 584960 6624
rect 579981 6566 584960 6568
rect 579981 6563 580047 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 214420 700708 214484 700772
rect 211660 700572 211724 700636
rect 215892 700436 215956 700500
rect 395292 700436 395356 700500
rect 213132 700300 213196 700364
rect 398604 700300 398668 700364
rect 397500 699816 397564 699820
rect 397500 699760 397514 699816
rect 397514 699760 397564 699816
rect 397500 699756 397564 699760
rect 170812 685944 170876 685948
rect 170812 685888 170862 685944
rect 170862 685888 170876 685944
rect 170812 685884 170876 685888
rect 350948 685944 351012 685948
rect 350948 685888 350998 685944
rect 350998 685888 351012 685944
rect 350948 685884 351012 685888
rect 530900 685944 530964 685948
rect 530900 685888 530950 685944
rect 530950 685888 530964 685944
rect 530900 685884 530964 685888
rect 38516 633388 38580 633452
rect 38332 608364 38396 608428
rect 38700 607412 38764 607476
rect 219204 607956 219268 608020
rect 357940 607412 358004 607476
rect 258086 599584 258150 599588
rect 258086 599528 258134 599584
rect 258134 599528 258150 599584
rect 258086 599524 258150 599528
rect 278486 599524 278550 599588
rect 435910 599584 435974 599588
rect 435910 599528 435914 599584
rect 435914 599528 435970 599584
rect 435970 599528 435974 599584
rect 435910 599524 435974 599528
rect 450860 599524 450924 599588
rect 451142 599524 451206 599588
rect 452148 599388 452212 599452
rect 61700 597484 61764 597548
rect 63172 597544 63236 597548
rect 63172 597488 63222 597544
rect 63222 597488 63236 597544
rect 63172 597484 63236 597488
rect 64276 597544 64340 597548
rect 64276 597488 64290 597544
rect 64290 597488 64340 597544
rect 64276 597484 64340 597488
rect 64644 597484 64708 597548
rect 66484 597484 66548 597548
rect 67588 597544 67652 597548
rect 67588 597488 67638 597544
rect 67638 597488 67652 597544
rect 67588 597484 67652 597488
rect 68324 597484 68388 597548
rect 69980 597484 70044 597548
rect 70716 597484 70780 597548
rect 73476 597484 73540 597548
rect 73660 597484 73724 597548
rect 74580 597484 74644 597548
rect 76052 597484 76116 597548
rect 78076 597544 78140 597548
rect 78076 597488 78090 597544
rect 78090 597488 78140 597544
rect 78076 597484 78140 597488
rect 78444 597484 78508 597548
rect 81020 597484 81084 597548
rect 83964 597484 84028 597548
rect 85988 597484 86052 597548
rect 88196 597544 88260 597548
rect 88196 597488 88246 597544
rect 88246 597488 88260 597544
rect 88196 597484 88260 597488
rect 93348 597484 93412 597548
rect 93532 597484 93596 597548
rect 122604 597484 122668 597548
rect 128492 597484 128556 597548
rect 131068 597544 131132 597548
rect 131068 597488 131082 597544
rect 131082 597488 131132 597544
rect 131068 597484 131132 597488
rect 133460 597484 133524 597548
rect 135852 597484 135916 597548
rect 141004 597484 141068 597548
rect 145972 597484 146036 597548
rect 235948 597544 236012 597548
rect 235948 597488 235998 597544
rect 235998 597488 236012 597544
rect 235948 597484 236012 597488
rect 237052 597484 237116 597548
rect 238156 597484 238220 597548
rect 243124 597544 243188 597548
rect 243124 597488 243138 597544
rect 243138 597488 243188 597544
rect 243124 597484 243188 597488
rect 244228 597544 244292 597548
rect 244228 597488 244278 597544
rect 244278 597488 244292 597544
rect 244228 597484 244292 597488
rect 245516 597544 245580 597548
rect 245516 597488 245530 597544
rect 245530 597488 245580 597544
rect 245516 597484 245580 597488
rect 246436 597544 246500 597548
rect 246436 597488 246486 597544
rect 246486 597488 246500 597544
rect 246436 597484 246500 597488
rect 248276 597484 248340 597548
rect 248644 597484 248708 597548
rect 250668 597484 250732 597548
rect 252324 597484 252388 597548
rect 253428 597544 253492 597548
rect 253428 597488 253478 597544
rect 253478 597488 253492 597544
rect 253428 597484 253492 597488
rect 254532 597544 254596 597548
rect 254532 597488 254582 597544
rect 254582 597488 254596 597544
rect 254532 597484 254596 597488
rect 255820 597484 255884 597548
rect 256924 597484 256988 597548
rect 261708 597484 261772 597548
rect 263548 597544 263612 597548
rect 263548 597488 263598 597544
rect 263598 597488 263612 597544
rect 263548 597484 263612 597488
rect 265940 597484 266004 597548
rect 268332 597484 268396 597548
rect 270908 597484 270972 597548
rect 276980 597484 277044 597548
rect 280844 597484 280908 597548
rect 283420 597484 283484 597548
rect 285996 597484 286060 597548
rect 290964 597484 291028 597548
rect 293356 597484 293420 597548
rect 416084 597484 416148 597548
rect 417188 597484 417252 597548
rect 418292 597484 418356 597548
rect 420500 597484 420564 597548
rect 421788 597484 421852 597548
rect 423076 597544 423140 597548
rect 423076 597488 423126 597544
rect 423126 597488 423140 597544
rect 423076 597484 423140 597488
rect 424180 597484 424244 597548
rect 425468 597484 425532 597548
rect 426572 597544 426636 597548
rect 426572 597488 426586 597544
rect 426586 597488 426636 597544
rect 426572 597484 426636 597488
rect 427676 597544 427740 597548
rect 427676 597488 427690 597544
rect 427690 597488 427740 597544
rect 427676 597484 427740 597488
rect 428596 597484 428660 597548
rect 430068 597484 430132 597548
rect 430620 597544 430684 597548
rect 430620 597488 430634 597544
rect 430634 597488 430684 597544
rect 430620 597484 430684 597488
rect 433748 597484 433812 597548
rect 434484 597544 434548 597548
rect 434484 597488 434534 597544
rect 434534 597488 434548 597544
rect 434484 597484 434548 597488
rect 435956 597484 436020 597548
rect 437060 597544 437124 597548
rect 437060 597488 437110 597544
rect 437110 597488 437124 597544
rect 437060 597484 437124 597488
rect 437980 597484 438044 597548
rect 439452 597484 439516 597548
rect 442764 597484 442828 597548
rect 443500 597484 443564 597548
rect 443868 597484 443932 597548
rect 445340 597484 445404 597548
rect 445892 597484 445956 597548
rect 448284 597484 448348 597548
rect 451044 597484 451108 597548
rect 58204 597348 58268 597412
rect 68692 597348 68756 597412
rect 71268 597408 71332 597412
rect 71268 597352 71318 597408
rect 71318 597352 71332 597408
rect 71268 597348 71332 597352
rect 72372 597348 72436 597412
rect 75868 597348 75932 597412
rect 76972 597348 77036 597412
rect 83780 597348 83844 597412
rect 39804 597212 39868 597276
rect 60596 597212 60660 597276
rect 81756 597212 81820 597276
rect 57100 597076 57164 597140
rect 59492 597076 59556 597140
rect 98132 597348 98196 597412
rect 108252 597348 108316 597412
rect 115980 597348 116044 597412
rect 120948 597348 121012 597412
rect 260972 597348 261036 597412
rect 262812 597348 262876 597412
rect 263916 597348 263980 597412
rect 267596 597348 267660 597412
rect 276060 597348 276124 597412
rect 300900 597348 300964 597412
rect 357572 597348 357636 597412
rect 456012 597484 456076 597548
rect 463556 597484 463620 597548
rect 465948 597484 466012 597548
rect 468156 597484 468220 597548
rect 473492 597484 473556 597548
rect 475884 597484 475948 597548
rect 478460 597484 478524 597548
rect 483428 597484 483492 597548
rect 486004 597484 486068 597548
rect 488580 597544 488644 597548
rect 488580 597488 488594 597544
rect 488594 597488 488644 597544
rect 488580 597484 488644 597488
rect 495940 597484 496004 597548
rect 498516 597484 498580 597548
rect 500908 597544 500972 597548
rect 500908 597488 500958 597544
rect 500958 597488 500972 597544
rect 500908 597484 500972 597488
rect 453252 597348 453316 597412
rect 86356 597212 86420 597276
rect 87644 597212 87708 597276
rect 95740 597212 95804 597276
rect 88748 597076 88812 597140
rect 89852 597076 89916 597140
rect 99052 597212 99116 597276
rect 113404 597212 113468 597276
rect 219020 597212 219084 597276
rect 273484 597212 273548 597276
rect 275692 597212 275756 597276
rect 298508 597212 298572 597276
rect 358860 597212 358924 597276
rect 460980 597212 461044 597276
rect 79364 596940 79428 597004
rect 80652 596940 80716 597004
rect 97028 597076 97092 597140
rect 125916 597076 125980 597140
rect 138428 597076 138492 597140
rect 271092 597076 271156 597140
rect 273300 597136 273364 597140
rect 273300 597080 273314 597136
rect 273314 597080 273364 597136
rect 273300 597076 273364 597080
rect 288204 597076 288268 597140
rect 357020 597076 357084 597140
rect 438532 597076 438596 597140
rect 440740 597076 440804 597140
rect 459140 597076 459204 597140
rect 111012 596940 111076 597004
rect 118556 597000 118620 597004
rect 118556 596944 118606 597000
rect 118606 596944 118620 597000
rect 118556 596940 118620 596944
rect 141924 596940 141988 597004
rect 325924 596940 325988 597004
rect 356652 596940 356716 597004
rect 441108 596940 441172 597004
rect 441660 597000 441724 597004
rect 441660 596944 441674 597000
rect 441674 596944 441724 597000
rect 441660 596940 441724 596944
rect 446260 596940 446324 597004
rect 447548 596940 447612 597004
rect 448652 596940 448716 597004
rect 454356 596940 454420 597004
rect 455644 596940 455708 597004
rect 480852 596940 480916 597004
rect 503300 596940 503364 597004
rect 82860 596864 82924 596868
rect 82860 596808 82874 596864
rect 82874 596808 82924 596864
rect 82860 596804 82924 596808
rect 103284 596804 103348 596868
rect 219940 596804 220004 596868
rect 238524 596804 238588 596868
rect 240548 596804 240612 596868
rect 241652 596804 241716 596868
rect 247540 596804 247604 596868
rect 250116 596804 250180 596868
rect 251404 596804 251468 596868
rect 265204 596804 265268 596868
rect 55996 596668 56060 596732
rect 100892 596668 100956 596732
rect 257844 596668 257908 596732
rect 259500 596728 259564 596732
rect 278084 596804 278148 596868
rect 311020 596804 311084 596868
rect 320956 596804 321020 596868
rect 323348 596804 323412 596868
rect 458404 596804 458468 596868
rect 505876 596804 505940 596868
rect 259500 596672 259550 596728
rect 259550 596672 259564 596728
rect 259500 596668 259564 596672
rect 268700 596668 268764 596732
rect 269804 596668 269868 596732
rect 313412 596668 313476 596732
rect 318564 596668 318628 596732
rect 419580 596728 419644 596732
rect 419580 596672 419594 596728
rect 419594 596672 419644 596728
rect 419580 596668 419644 596672
rect 428228 596668 428292 596732
rect 431172 596668 431236 596732
rect 431908 596728 431972 596732
rect 431908 596672 431958 596728
rect 431958 596672 431972 596728
rect 431908 596668 431972 596672
rect 433380 596728 433444 596732
rect 433380 596672 433430 596728
rect 433430 596672 433444 596728
rect 433380 596668 433444 596672
rect 458036 596668 458100 596732
rect 493364 596668 493428 596732
rect 92244 596532 92308 596596
rect 94452 596532 94516 596596
rect 106044 596532 106108 596596
rect 216260 596532 216324 596596
rect 256004 596532 256068 596596
rect 260604 596532 260668 596596
rect 279188 596532 279252 596596
rect 315804 596532 315868 596596
rect 83596 596396 83660 596460
rect 91140 596456 91204 596460
rect 91140 596400 91154 596456
rect 91154 596400 91204 596456
rect 91140 596396 91204 596400
rect 96108 596396 96172 596460
rect 98500 596396 98564 596460
rect 266308 596456 266372 596460
rect 266308 596400 266358 596456
rect 266358 596400 266372 596456
rect 266308 596396 266372 596400
rect 272196 596396 272260 596460
rect 306052 596456 306116 596460
rect 306052 596400 306102 596456
rect 306102 596400 306116 596456
rect 306052 596396 306116 596400
rect 308628 596396 308692 596460
rect 453620 596532 453684 596596
rect 450860 596396 450924 596460
rect 90956 596320 91020 596324
rect 90956 596264 91006 596320
rect 91006 596264 91020 596320
rect 90956 596260 91020 596264
rect 210740 596260 210804 596324
rect 253612 596260 253676 596324
rect 274404 596260 274468 596324
rect 295932 596260 295996 596324
rect 303476 596320 303540 596324
rect 303476 596264 303526 596320
rect 303526 596264 303540 596320
rect 303476 596260 303540 596264
rect 449756 596260 449820 596324
rect 456932 596260 456996 596324
rect 470364 596260 470428 596324
rect 489684 596260 489748 596324
rect 399340 594492 399404 594556
rect 215156 594084 215220 594148
rect 217732 593948 217796 594012
rect 358124 592588 358188 592652
rect 212396 571916 212460 571980
rect 218652 570692 218716 570756
rect 216444 570556 216508 570620
rect 217916 567156 217980 567220
rect 210924 566476 210988 566540
rect 212580 566340 212644 566404
rect 170812 565856 170876 565860
rect 170812 565800 170862 565856
rect 170862 565800 170876 565856
rect 170812 565796 170876 565800
rect 350948 565796 351012 565860
rect 530900 565856 530964 565860
rect 530900 565800 530950 565856
rect 530950 565800 530964 565856
rect 530900 565796 530964 565800
rect 203380 565388 203444 565452
rect 206140 565252 206204 565316
rect 206324 565116 206388 565180
rect 208716 564980 208780 565044
rect 219756 563620 219820 563684
rect 38516 514040 38580 514044
rect 38516 513984 38530 514040
rect 38530 513984 38580 514040
rect 38516 513980 38580 513984
rect 397132 513708 397196 513772
rect 38332 488276 38396 488340
rect 217916 488276 217980 488340
rect 38884 487460 38948 487524
rect 397316 487324 397380 487388
rect 217916 487188 217980 487252
rect 359412 487188 359476 487252
rect 56054 479632 56118 479636
rect 56054 479576 56102 479632
rect 56102 479576 56118 479632
rect 56054 479572 56118 479576
rect 236054 479572 236118 479636
rect 217180 478892 217244 478956
rect 72372 478680 72436 478684
rect 72372 478624 72386 478680
rect 72386 478624 72436 478680
rect 72372 478620 72436 478624
rect 74580 478680 74644 478684
rect 74580 478624 74630 478680
rect 74630 478624 74644 478680
rect 74580 478620 74644 478624
rect 73476 478484 73540 478548
rect 76972 478544 77036 478548
rect 76972 478488 76986 478544
rect 76986 478488 77036 478544
rect 76972 478484 77036 478488
rect 75868 478408 75932 478412
rect 75868 478352 75882 478408
rect 75882 478352 75932 478408
rect 75868 478348 75932 478352
rect 428596 478408 428660 478412
rect 428596 478352 428610 478408
rect 428610 478352 428660 478408
rect 428596 478348 428660 478352
rect 430068 478408 430132 478412
rect 430068 478352 430118 478408
rect 430118 478352 430132 478408
rect 430068 478348 430132 478352
rect 79548 478272 79612 478276
rect 79548 478216 79562 478272
rect 79562 478216 79612 478272
rect 79548 478212 79612 478216
rect 431356 478272 431420 478276
rect 431356 478216 431370 478272
rect 431370 478216 431420 478272
rect 431356 478212 431420 478216
rect 432460 478272 432524 478276
rect 432460 478216 432510 478272
rect 432510 478216 432524 478272
rect 432460 478212 432524 478216
rect 80652 478136 80716 478140
rect 80652 478080 80666 478136
rect 80666 478080 80716 478136
rect 80652 478076 80716 478080
rect 86356 477592 86420 477596
rect 86356 477536 86370 477592
rect 86370 477536 86420 477592
rect 86356 477532 86420 477536
rect 39804 477396 39868 477460
rect 60596 477396 60660 477460
rect 63172 477456 63236 477460
rect 63172 477400 63222 477456
rect 63222 477400 63236 477456
rect 63172 477396 63236 477400
rect 64276 477456 64340 477460
rect 64276 477400 64290 477456
rect 64290 477400 64340 477456
rect 64276 477396 64340 477400
rect 65380 477396 65444 477460
rect 66484 477456 66548 477460
rect 66484 477400 66534 477456
rect 66534 477400 66548 477456
rect 66484 477396 66548 477400
rect 67588 477456 67652 477460
rect 67588 477400 67638 477456
rect 67638 477400 67652 477456
rect 67588 477396 67652 477400
rect 68692 477456 68756 477460
rect 68692 477400 68742 477456
rect 68742 477400 68756 477456
rect 68692 477396 68756 477400
rect 70164 477456 70228 477460
rect 70164 477400 70214 477456
rect 70214 477400 70228 477456
rect 70164 477396 70228 477400
rect 71268 477396 71332 477460
rect 78076 477456 78140 477460
rect 78076 477400 78126 477456
rect 78126 477400 78140 477456
rect 78076 477396 78140 477400
rect 81020 477396 81084 477460
rect 81756 477456 81820 477460
rect 81756 477400 81806 477456
rect 81806 477400 81820 477456
rect 81756 477396 81820 477400
rect 82860 477456 82924 477460
rect 82860 477400 82874 477456
rect 82874 477400 82924 477456
rect 82860 477396 82924 477400
rect 83596 477396 83660 477460
rect 85252 477456 85316 477460
rect 85252 477400 85302 477456
rect 85302 477400 85316 477456
rect 85252 477396 85316 477400
rect 85988 477396 86052 477460
rect 87644 477456 87708 477460
rect 87644 477400 87658 477456
rect 87658 477400 87708 477456
rect 87644 477396 87708 477400
rect 88196 477456 88260 477460
rect 88196 477400 88246 477456
rect 88246 477400 88260 477456
rect 88196 477396 88260 477400
rect 88748 477456 88812 477460
rect 88748 477400 88762 477456
rect 88762 477400 88812 477456
rect 88748 477396 88812 477400
rect 89852 477396 89916 477460
rect 91140 477456 91204 477460
rect 91140 477400 91190 477456
rect 91190 477400 91204 477456
rect 91140 477396 91204 477400
rect 92244 477456 92308 477460
rect 92244 477400 92258 477456
rect 92258 477400 92308 477456
rect 92244 477396 92308 477400
rect 93348 477396 93412 477460
rect 94452 477456 94516 477460
rect 94452 477400 94466 477456
rect 94466 477400 94516 477456
rect 94452 477396 94516 477400
rect 95740 477456 95804 477460
rect 95740 477400 95790 477456
rect 95790 477400 95804 477456
rect 95740 477396 95804 477400
rect 97028 477456 97092 477460
rect 97028 477400 97042 477456
rect 97042 477400 97092 477456
rect 97028 477396 97092 477400
rect 99052 477396 99116 477460
rect 59492 477320 59556 477324
rect 59492 477264 59506 477320
rect 59506 477264 59556 477320
rect 59492 477260 59556 477264
rect 61700 477260 61764 477324
rect 239628 477396 239692 477460
rect 243124 477456 243188 477460
rect 243124 477400 243174 477456
rect 243174 477400 243188 477456
rect 243124 477396 243188 477400
rect 244228 477456 244292 477460
rect 244228 477400 244278 477456
rect 244278 477400 244292 477456
rect 244228 477396 244292 477400
rect 245516 477456 245580 477460
rect 245516 477400 245530 477456
rect 245530 477400 245580 477456
rect 245516 477396 245580 477400
rect 246436 477396 246500 477460
rect 247540 477396 247604 477460
rect 248644 477456 248708 477460
rect 248644 477400 248658 477456
rect 248658 477400 248708 477456
rect 248644 477396 248708 477400
rect 250116 477456 250180 477460
rect 250116 477400 250130 477456
rect 250130 477400 250180 477456
rect 250116 477396 250180 477400
rect 251220 477456 251284 477460
rect 251220 477400 251270 477456
rect 251270 477400 251284 477456
rect 251220 477396 251284 477400
rect 252324 477456 252388 477460
rect 252324 477400 252374 477456
rect 252374 477400 252388 477456
rect 252324 477396 252388 477400
rect 253428 477456 253492 477460
rect 253428 477400 253442 477456
rect 253442 477400 253492 477456
rect 253428 477396 253492 477400
rect 254532 477456 254596 477460
rect 254532 477400 254546 477456
rect 254546 477400 254596 477456
rect 254532 477396 254596 477400
rect 255820 477396 255884 477460
rect 256924 477456 256988 477460
rect 256924 477400 256974 477456
rect 256974 477400 256988 477456
rect 256924 477396 256988 477400
rect 260788 477456 260852 477460
rect 260788 477400 260838 477456
rect 260838 477400 260852 477456
rect 260788 477396 260852 477400
rect 266308 477456 266372 477460
rect 266308 477400 266358 477456
rect 266358 477400 266372 477456
rect 266308 477396 266372 477400
rect 269804 477396 269868 477460
rect 279188 477396 279252 477460
rect 416084 477396 416148 477460
rect 417188 477396 417252 477460
rect 418292 477396 418356 477460
rect 420500 477396 420564 477460
rect 421788 477396 421852 477460
rect 423076 477456 423140 477460
rect 423076 477400 423126 477456
rect 423126 477400 423140 477456
rect 423076 477396 423140 477400
rect 424180 477456 424244 477460
rect 424180 477400 424194 477456
rect 424194 477400 424244 477456
rect 424180 477396 424244 477400
rect 425468 477456 425532 477460
rect 425468 477400 425518 477456
rect 425518 477400 425532 477456
rect 425468 477396 425532 477400
rect 426572 477456 426636 477460
rect 426572 477400 426622 477456
rect 426622 477400 426636 477456
rect 426572 477396 426636 477400
rect 427676 477456 427740 477460
rect 427676 477400 427726 477456
rect 427726 477400 427740 477456
rect 427676 477396 427740 477400
rect 433380 477456 433444 477460
rect 433380 477400 433430 477456
rect 433430 477400 433444 477456
rect 433380 477396 433444 477400
rect 434484 477456 434548 477460
rect 434484 477400 434534 477456
rect 434534 477400 434548 477456
rect 434484 477396 434548 477400
rect 435772 477456 435836 477460
rect 435772 477400 435786 477456
rect 435786 477400 435836 477456
rect 435772 477396 435836 477400
rect 437060 477396 437124 477460
rect 438164 477456 438228 477460
rect 438164 477400 438178 477456
rect 438178 477400 438228 477456
rect 438164 477396 438228 477400
rect 443868 477396 443932 477460
rect 447548 477396 447612 477460
rect 449756 477396 449820 477460
rect 453252 477396 453316 477460
rect 237052 477260 237116 477324
rect 258212 477260 258276 477324
rect 261708 477260 261772 477324
rect 263916 477260 263980 477324
rect 272196 477260 272260 477324
rect 276980 477260 277044 477324
rect 278084 477260 278148 477324
rect 460980 477260 461044 477324
rect 241652 477124 241716 477188
rect 274404 477124 274468 477188
rect 275692 477124 275756 477188
rect 311020 477124 311084 477188
rect 435956 477124 436020 477188
rect 439452 477124 439516 477188
rect 445340 477124 445404 477188
rect 446260 477124 446324 477188
rect 448652 477124 448716 477188
rect 452148 477124 452212 477188
rect 459140 477124 459204 477188
rect 463556 477124 463620 477188
rect 60596 476988 60660 477052
rect 240548 476988 240612 477052
rect 265204 476988 265268 477052
rect 271276 476988 271340 477052
rect 278452 476988 278516 477052
rect 285996 476988 286060 477052
rect 323348 476988 323412 477052
rect 325924 476988 325988 477052
rect 438532 476988 438596 477052
rect 440740 476988 440804 477052
rect 453620 476988 453684 477052
rect 454356 476988 454420 477052
rect 456932 476988 456996 477052
rect 58204 476912 58268 476916
rect 58204 476856 58218 476912
rect 58218 476856 58268 476912
rect 58204 476852 58268 476856
rect 238156 476852 238220 476916
rect 256188 476852 256252 476916
rect 262812 476852 262876 476916
rect 270908 476852 270972 476916
rect 273300 476912 273364 476916
rect 273300 476856 273314 476912
rect 273314 476856 273364 476912
rect 273300 476852 273364 476856
rect 320956 476852 321020 476916
rect 441108 476852 441172 476916
rect 441660 476912 441724 476916
rect 441660 476856 441674 476912
rect 441674 476856 441724 476912
rect 441660 476852 441724 476856
rect 455644 476852 455708 476916
rect 458036 476852 458100 476916
rect 483428 476852 483492 476916
rect 57100 476716 57164 476780
rect 267596 476716 267660 476780
rect 288204 476716 288268 476780
rect 300900 476716 300964 476780
rect 315804 476716 315868 476780
rect 318564 476716 318628 476780
rect 456012 476716 456076 476780
rect 490972 476716 491036 476780
rect 498516 476716 498580 476780
rect 83964 476640 84028 476644
rect 83964 476584 84014 476640
rect 84014 476584 84028 476640
rect 83964 476580 84028 476584
rect 90956 476504 91020 476508
rect 90956 476448 91006 476504
rect 91006 476448 91020 476504
rect 90956 476444 91020 476448
rect 93532 476444 93596 476508
rect 99052 476444 99116 476508
rect 79548 476308 79612 476372
rect 98132 476308 98196 476372
rect 259500 476580 259564 476644
rect 268700 476580 268764 476644
rect 308628 476580 308692 476644
rect 313412 476580 313476 476644
rect 260788 476444 260852 476508
rect 290964 476444 291028 476508
rect 306052 476504 306116 476508
rect 306052 476448 306102 476504
rect 306102 476448 306116 476504
rect 306052 476444 306116 476448
rect 419580 476504 419644 476508
rect 419580 476448 419594 476504
rect 419594 476448 419644 476504
rect 419580 476444 419644 476448
rect 433748 476444 433812 476508
rect 442764 476444 442828 476508
rect 443500 476444 443564 476508
rect 451044 476444 451108 476508
rect 475884 476444 475948 476508
rect 478460 476444 478524 476508
rect 298508 476308 298572 476372
rect 303476 476368 303540 476372
rect 303476 476312 303526 476368
rect 303526 476312 303540 476368
rect 303476 476308 303540 476312
rect 458404 476308 458468 476372
rect 503300 476308 503364 476372
rect 68324 476172 68388 476236
rect 70716 476172 70780 476236
rect 73660 476172 73724 476236
rect 76052 476172 76116 476236
rect 78444 476172 78508 476236
rect 96108 476172 96172 476236
rect 98500 476172 98564 476236
rect 100892 476172 100956 476236
rect 103652 476172 103716 476236
rect 106044 476172 106108 476236
rect 108252 476172 108316 476236
rect 111012 476172 111076 476236
rect 113404 476172 113468 476236
rect 115980 476172 116044 476236
rect 118556 476232 118620 476236
rect 118556 476176 118606 476232
rect 118606 476176 118620 476232
rect 118556 476172 118620 476176
rect 120948 476172 121012 476236
rect 123524 476172 123588 476236
rect 125916 476172 125980 476236
rect 128492 476172 128556 476236
rect 131068 476232 131132 476236
rect 131068 476176 131082 476232
rect 131082 476176 131132 476232
rect 131068 476172 131132 476176
rect 133460 476172 133524 476236
rect 135852 476172 135916 476236
rect 138428 476172 138492 476236
rect 141004 476172 141068 476236
rect 143396 476232 143460 476236
rect 143396 476176 143446 476232
rect 143446 476176 143460 476232
rect 143396 476172 143460 476176
rect 145972 476172 146036 476236
rect 248276 476172 248340 476236
rect 250668 476172 250732 476236
rect 253612 476172 253676 476236
rect 258396 476172 258460 476236
rect 260972 476172 261036 476236
rect 263548 476232 263612 476236
rect 263548 476176 263598 476232
rect 263598 476176 263612 476232
rect 263548 476172 263612 476176
rect 265940 476172 266004 476236
rect 268332 476172 268396 476236
rect 273484 476172 273548 476236
rect 276060 476232 276124 476236
rect 276060 476176 276074 476232
rect 276074 476176 276124 476232
rect 276060 476172 276124 476176
rect 280844 476172 280908 476236
rect 283420 476172 283484 476236
rect 293356 476172 293420 476236
rect 295932 476172 295996 476236
rect 428228 476172 428292 476236
rect 430620 476232 430684 476236
rect 430620 476176 430634 476232
rect 430634 476176 430684 476232
rect 430620 476172 430684 476176
rect 445892 476172 445956 476236
rect 448284 476172 448348 476236
rect 450860 476172 450924 476236
rect 465948 476172 466012 476236
rect 468156 476172 468220 476236
rect 470916 476172 470980 476236
rect 473492 476172 473556 476236
rect 480852 476172 480916 476236
rect 486004 476172 486068 476236
rect 488580 476232 488644 476236
rect 488580 476176 488594 476232
rect 488594 476176 488644 476232
rect 488580 476172 488644 476176
rect 493364 476172 493428 476236
rect 495940 476172 496004 476236
rect 500908 476232 500972 476236
rect 500908 476176 500958 476232
rect 500958 476176 500972 476232
rect 500908 476172 500972 476176
rect 505876 476172 505940 476236
rect 217732 474676 217796 474740
rect 218836 474676 218900 474740
rect 399524 474540 399588 474604
rect 216076 461484 216140 461548
rect 212212 460124 212276 460188
rect 397316 446388 397380 446452
rect 530900 446388 530964 446452
rect 170812 445768 170876 445772
rect 170812 445712 170862 445768
rect 170862 445712 170876 445768
rect 170812 445708 170876 445712
rect 350948 445708 351012 445772
rect 214788 445164 214852 445228
rect 214604 445028 214668 445092
rect 216812 444892 216876 444956
rect 398788 444212 398852 444276
rect 216628 443532 216692 443596
rect 397132 394572 397196 394636
rect 217732 393892 217796 393956
rect 217180 393756 217244 393820
rect 217364 369956 217428 370020
rect 216812 369880 216876 369884
rect 216812 369824 216862 369880
rect 216862 369824 216876 369880
rect 216812 369820 216876 369824
rect 217548 368324 217612 368388
rect 217916 368324 217980 368388
rect 397316 368324 397380 368388
rect 219204 359892 219268 359956
rect 217732 359620 217796 359684
rect 357572 359484 357636 359548
rect 450860 359484 450924 359548
rect 451142 359484 451206 359548
rect 218836 359348 218900 359412
rect 358860 359348 358924 359412
rect 216260 358668 216324 358732
rect 325924 358668 325988 358732
rect 235948 358592 236012 358596
rect 235948 358536 235998 358592
rect 235998 358536 236012 358592
rect 235948 358532 236012 358536
rect 210740 358396 210804 358460
rect 60596 358124 60660 358188
rect 64276 358184 64340 358188
rect 64276 358128 64326 358184
rect 64326 358128 64340 358184
rect 64276 358124 64340 358128
rect 219020 358124 219084 358188
rect 276060 358184 276124 358188
rect 276060 358128 276074 358184
rect 276074 358128 276124 358184
rect 276060 358124 276124 358128
rect 300900 358184 300964 358188
rect 300900 358128 300914 358184
rect 300914 358128 300964 358184
rect 300900 358124 300964 358128
rect 416084 358184 416148 358188
rect 416084 358128 416098 358184
rect 416098 358128 416148 358184
rect 416084 358124 416148 358128
rect 488580 358184 488644 358188
rect 488580 358128 488594 358184
rect 488594 358128 488644 358184
rect 488580 358124 488644 358128
rect 55996 357308 56060 357372
rect 58204 357308 58268 357372
rect 59676 357308 59740 357372
rect 61884 357308 61948 357372
rect 63172 357308 63236 357372
rect 66484 357308 66548 357372
rect 68692 357308 68756 357372
rect 70164 357308 70228 357372
rect 71268 357308 71332 357372
rect 72372 357308 72436 357372
rect 73476 357308 73540 357372
rect 74580 357308 74644 357372
rect 76972 357308 77036 357372
rect 78444 357308 78508 357372
rect 79548 357308 79612 357372
rect 81020 357308 81084 357372
rect 85988 357308 86052 357372
rect 88196 357368 88260 357372
rect 88196 357312 88246 357368
rect 88246 357312 88260 357368
rect 88196 357308 88260 357312
rect 90956 357368 91020 357372
rect 90956 357312 91006 357368
rect 91006 357312 91020 357368
rect 90956 357308 91020 357312
rect 93532 357308 93596 357372
rect 95924 357308 95988 357372
rect 98500 357308 98564 357372
rect 100892 357308 100956 357372
rect 106044 357308 106108 357372
rect 243124 357308 243188 357372
rect 248276 357308 248340 357372
rect 248644 357368 248708 357372
rect 248644 357312 248694 357368
rect 248694 357312 248708 357368
rect 248644 357308 248708 357312
rect 250668 357308 250732 357372
rect 251220 357368 251284 357372
rect 251220 357312 251270 357368
rect 251270 357312 251284 357368
rect 251220 357308 251284 357312
rect 253612 357308 253676 357372
rect 254532 357368 254596 357372
rect 254532 357312 254582 357368
rect 254582 357312 254596 357368
rect 254532 357308 254596 357312
rect 256004 357308 256068 357372
rect 257108 357308 257172 357372
rect 258396 357308 258460 357372
rect 260972 357308 261036 357372
rect 262076 357368 262140 357372
rect 262076 357312 262126 357368
rect 262126 357312 262140 357368
rect 262076 357308 262140 357312
rect 262812 357368 262876 357372
rect 262812 357312 262826 357368
rect 262826 357312 262876 357368
rect 262812 357308 262876 357312
rect 263548 357308 263612 357372
rect 263916 357368 263980 357372
rect 263916 357312 263966 357368
rect 263966 357312 263980 357368
rect 263916 357308 263980 357312
rect 265756 357368 265820 357372
rect 265756 357312 265770 357368
rect 265770 357312 265820 357368
rect 265756 357308 265820 357312
rect 266308 357308 266372 357372
rect 267596 357368 267660 357372
rect 267596 357312 267610 357368
rect 267610 357312 267660 357368
rect 267596 357308 267660 357312
rect 268332 357308 268396 357372
rect 268516 357368 268580 357372
rect 268516 357312 268566 357368
rect 268566 357312 268580 357368
rect 268516 357308 268580 357312
rect 269804 357368 269868 357372
rect 269804 357312 269818 357368
rect 269818 357312 269868 357368
rect 269804 357308 269868 357312
rect 270908 357308 270972 357372
rect 271092 357368 271156 357372
rect 271092 357312 271142 357368
rect 271142 357312 271156 357368
rect 271092 357308 271156 357312
rect 272196 357368 272260 357372
rect 272196 357312 272210 357368
rect 272210 357312 272260 357368
rect 272196 357308 272260 357312
rect 273300 357368 273364 357372
rect 273300 357312 273350 357368
rect 273350 357312 273364 357368
rect 273300 357308 273364 357312
rect 274404 357308 274468 357372
rect 275876 357368 275940 357372
rect 275876 357312 275926 357368
rect 275926 357312 275940 357368
rect 275876 357308 275940 357312
rect 276980 357368 277044 357372
rect 276980 357312 277030 357368
rect 277030 357312 277044 357368
rect 276980 357308 277044 357312
rect 283420 357308 283484 357372
rect 285996 357308 286060 357372
rect 288204 357308 288268 357372
rect 290964 357308 291028 357372
rect 293356 357308 293420 357372
rect 295932 357308 295996 357372
rect 298508 357308 298572 357372
rect 303476 357308 303540 357372
rect 305868 357308 305932 357372
rect 308076 357308 308140 357372
rect 311020 357308 311084 357372
rect 313412 357308 313476 357372
rect 315620 357308 315684 357372
rect 318380 357308 318444 357372
rect 320956 357308 321020 357372
rect 417188 357308 417252 357372
rect 423076 357368 423140 357372
rect 423076 357312 423126 357368
rect 423126 357312 423140 357368
rect 423076 357308 423140 357312
rect 424548 357308 424612 357372
rect 425468 357368 425532 357372
rect 425468 357312 425482 357368
rect 425482 357312 425532 357368
rect 425468 357308 425532 357312
rect 426572 357308 426636 357372
rect 427676 357368 427740 357372
rect 427676 357312 427690 357368
rect 427690 357312 427740 357368
rect 427676 357308 427740 357312
rect 428228 357308 428292 357372
rect 428596 357368 428660 357372
rect 428596 357312 428610 357368
rect 428610 357312 428660 357368
rect 428596 357308 428660 357312
rect 430068 357368 430132 357372
rect 430068 357312 430082 357368
rect 430082 357312 430132 357368
rect 430068 357308 430132 357312
rect 430620 357368 430684 357372
rect 430620 357312 430634 357368
rect 430634 357312 430684 357368
rect 430620 357308 430684 357312
rect 431908 357368 431972 357372
rect 431908 357312 431958 357368
rect 431958 357312 431972 357368
rect 431908 357308 431972 357312
rect 433564 357308 433628 357372
rect 435956 357308 436020 357372
rect 437060 357308 437124 357372
rect 438532 357308 438596 357372
rect 440924 357308 440988 357372
rect 445892 357368 445956 357372
rect 445892 357312 445906 357368
rect 445906 357312 445956 357368
rect 57100 357172 57164 357236
rect 70716 357172 70780 357236
rect 73292 357172 73356 357236
rect 75868 357172 75932 357236
rect 78260 357172 78324 357236
rect 80652 357172 80716 357236
rect 238340 357172 238404 357236
rect 418108 357172 418172 357236
rect 431172 357172 431236 357236
rect 433380 357232 433444 357236
rect 433380 357176 433430 357232
rect 433430 357176 433444 357232
rect 433380 357172 433444 357176
rect 434668 357232 434732 357236
rect 434668 357176 434682 357232
rect 434682 357176 434732 357232
rect 434668 357172 434732 357176
rect 435772 357172 435836 357236
rect 438348 357232 438412 357236
rect 438348 357176 438398 357232
rect 438398 357176 438412 357232
rect 438348 357172 438412 357176
rect 438900 357172 438964 357236
rect 439452 357172 439516 357236
rect 445892 357308 445956 357312
rect 448284 357308 448348 357372
rect 451044 357308 451108 357372
rect 452148 357308 452212 357372
rect 453620 357308 453684 357372
rect 455828 357308 455892 357372
rect 458404 357308 458468 357372
rect 463556 357308 463620 357372
rect 465948 357308 466012 357372
rect 468156 357308 468220 357372
rect 473308 357308 473372 357372
rect 478460 357308 478524 357372
rect 486004 357308 486068 357372
rect 498516 357308 498580 357372
rect 443500 357172 443564 357236
rect 458036 357172 458100 357236
rect 459140 357172 459204 357236
rect 68324 357036 68388 357100
rect 238892 357036 238956 357100
rect 419580 357036 419644 357100
rect 244596 356900 244660 356964
rect 419948 356900 420012 356964
rect 83596 356628 83660 356692
rect 241836 356764 241900 356828
rect 421788 356764 421852 356828
rect 245516 356688 245580 356692
rect 245516 356632 245566 356688
rect 245566 356632 245580 356688
rect 245516 356628 245580 356632
rect 250116 356688 250180 356692
rect 250116 356632 250130 356688
rect 250130 356632 250180 356688
rect 250116 356628 250180 356632
rect 252324 356688 252388 356692
rect 252324 356632 252338 356688
rect 252338 356632 252388 356688
rect 252324 356628 252388 356632
rect 255820 356688 255884 356692
rect 255820 356632 255834 356688
rect 255834 356632 255884 356688
rect 255820 356628 255884 356632
rect 258396 356628 258460 356692
rect 259500 356628 259564 356692
rect 278084 356628 278148 356692
rect 247540 356492 247604 356556
rect 253428 356552 253492 356556
rect 253428 356496 253442 356552
rect 253442 356496 253492 356552
rect 253428 356492 253492 356496
rect 265940 356492 266004 356556
rect 76052 356356 76116 356420
rect 246620 356356 246684 356420
rect 260604 356356 260668 356420
rect 279188 356492 279252 356556
rect 440740 356492 440804 356556
rect 447548 357036 447612 357100
rect 450860 357036 450924 357100
rect 454356 357036 454420 357100
rect 480668 357036 480732 357100
rect 453252 356900 453316 356964
rect 455644 356900 455708 356964
rect 448468 356824 448532 356828
rect 448468 356768 448518 356824
rect 448518 356768 448532 356824
rect 448468 356764 448532 356768
rect 456932 356764 456996 356828
rect 503300 356764 503364 356828
rect 446260 356628 446324 356692
rect 442028 356492 442092 356556
rect 443868 356492 443932 356556
rect 449756 356492 449820 356556
rect 483428 356492 483492 356556
rect 438900 356356 438964 356420
rect 442764 356356 442828 356420
rect 444788 356356 444852 356420
rect 475884 356356 475948 356420
rect 500908 356416 500972 356420
rect 500908 356360 500958 356416
rect 500958 356360 500972 356416
rect 500908 356356 500972 356360
rect 237236 356220 237300 356284
rect 470916 356220 470980 356284
rect 489684 356220 489748 356284
rect 495572 356220 495636 356284
rect 64644 356084 64708 356148
rect 67588 356084 67652 356148
rect 103284 356084 103348 356148
rect 240916 356084 240980 356148
rect 273484 356084 273548 356148
rect 278452 356084 278516 356148
rect 280844 356084 280908 356148
rect 323348 356084 323412 356148
rect 460980 356144 461044 356148
rect 460980 356088 460994 356144
rect 460994 356088 461044 356144
rect 460980 356084 461044 356088
rect 493364 356084 493428 356148
rect 505508 356084 505572 356148
rect 215156 355404 215220 355468
rect 215892 355268 215956 355332
rect 397500 352548 397564 352612
rect 399524 351188 399588 351252
rect 395292 351052 395356 351116
rect 398604 349692 398668 349756
rect 399340 348332 399404 348396
rect 211660 342892 211724 342956
rect 217364 342892 217428 342956
rect 213132 337316 213196 337380
rect 214420 327660 214484 327724
rect 38700 324940 38764 325004
rect 398788 311068 398852 311132
rect 38884 304132 38948 304196
rect 357020 298692 357084 298756
rect 356652 297332 356716 297396
rect 357940 294476 358004 294540
rect 206324 293524 206388 293588
rect 206140 293388 206204 293452
rect 203380 293252 203444 293316
rect 359412 293116 359476 293180
rect 219940 289036 220004 289100
rect 214604 287812 214668 287876
rect 214788 287676 214852 287740
rect 208716 282780 208780 282844
rect 210924 282780 210988 282844
rect 212212 282780 212276 282844
rect 216076 282780 216140 282844
rect 216444 282780 216508 282844
rect 216628 282780 216692 282844
rect 218652 282780 218716 282844
rect 219756 282780 219820 282844
rect 212396 282644 212460 282708
rect 212580 282644 212644 282708
rect 217548 282508 217612 282572
rect 358124 282236 358188 282300
rect 123708 279516 123772 279580
rect 123892 279244 123956 279308
rect 123708 31724 123772 31788
rect 123892 7516 123956 7580
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 24114 493774 24734 529218
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 169774 24734 205218
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 24114 25774 24734 61218
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 685244 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 685244 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 685244 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 685244 49574 698058
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 685244 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 685244 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 685244 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 685244 85574 698058
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 685244 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 685244 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 685244 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 685244 121574 698058
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 685244 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 685244 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 685244 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 685244 157574 698058
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 170811 685948 170877 685949
rect 170811 685884 170812 685948
rect 170876 685884 170877 685948
rect 170811 685883 170877 685884
rect 170814 683770 170874 685883
rect 170814 683710 170900 683770
rect 170840 683202 170900 683710
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 40272 655174 40620 655206
rect 40272 654938 40328 655174
rect 40564 654938 40620 655174
rect 40272 654854 40620 654938
rect 40272 654618 40328 654854
rect 40564 654618 40620 654854
rect 40272 654586 40620 654618
rect 176000 655174 176348 655206
rect 176000 654938 176056 655174
rect 176292 654938 176348 655174
rect 176000 654854 176348 654938
rect 176000 654618 176056 654854
rect 176292 654618 176348 654854
rect 176000 654586 176348 654618
rect 40952 651454 41300 651486
rect 40952 651218 41008 651454
rect 41244 651218 41300 651454
rect 40952 651134 41300 651218
rect 40952 650898 41008 651134
rect 41244 650898 41300 651134
rect 40952 650866 41300 650898
rect 175320 651454 175668 651486
rect 175320 651218 175376 651454
rect 175612 651218 175668 651454
rect 175320 651134 175668 651218
rect 175320 650898 175376 651134
rect 175612 650898 175668 651134
rect 175320 650866 175668 650898
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 605494 28454 640938
rect 38515 633452 38581 633453
rect 38515 633388 38516 633452
rect 38580 633388 38581 633452
rect 38515 633387 38581 633388
rect 38331 608428 38397 608429
rect 38331 608364 38332 608428
rect 38396 608364 38397 608428
rect 38331 608363 38397 608364
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 38334 488341 38394 608363
rect 38518 514045 38578 633387
rect 40272 619174 40620 619206
rect 40272 618938 40328 619174
rect 40564 618938 40620 619174
rect 40272 618854 40620 618938
rect 40272 618618 40328 618854
rect 40564 618618 40620 618854
rect 40272 618586 40620 618618
rect 176000 619174 176348 619206
rect 176000 618938 176056 619174
rect 176292 618938 176348 619174
rect 176000 618854 176348 618938
rect 176000 618618 176056 618854
rect 176292 618618 176348 618854
rect 176000 618586 176348 618618
rect 40952 615454 41300 615486
rect 40952 615218 41008 615454
rect 41244 615218 41300 615454
rect 40952 615134 41300 615218
rect 40952 614898 41008 615134
rect 41244 614898 41300 615134
rect 40952 614866 41300 614898
rect 175320 615454 175668 615486
rect 175320 615218 175376 615454
rect 175612 615218 175668 615454
rect 175320 615134 175668 615218
rect 175320 614898 175376 615134
rect 175612 614898 175668 615134
rect 175320 614866 175668 614898
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 38699 607476 38765 607477
rect 38699 607412 38700 607476
rect 38764 607412 38765 607476
rect 38699 607411 38765 607412
rect 38515 514044 38581 514045
rect 38515 513980 38516 514044
rect 38580 513980 38581 514044
rect 38515 513979 38581 513980
rect 38331 488340 38397 488341
rect 38331 488276 38332 488340
rect 38396 488276 38397 488340
rect 38331 488275 38397 488276
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 327454 38414 358064
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 38702 325005 38762 607411
rect 56056 599450 56116 600100
rect 57144 599450 57204 600100
rect 58232 599450 58292 600100
rect 59592 599450 59652 600100
rect 55998 599390 56116 599450
rect 57102 599390 57204 599450
rect 58206 599390 58292 599450
rect 59494 599390 59652 599450
rect 60544 599450 60604 600100
rect 61768 599450 61828 600100
rect 60544 599390 60658 599450
rect 39803 597276 39869 597277
rect 39803 597212 39804 597276
rect 39868 597212 39869 597276
rect 39803 597211 39869 597212
rect 38883 487524 38949 487525
rect 38883 487460 38884 487524
rect 38948 487460 38949 487524
rect 38883 487459 38949 487460
rect 38699 325004 38765 325005
rect 38699 324940 38700 325004
rect 38764 324940 38765 325004
rect 38699 324939 38765 324940
rect 38886 304197 38946 487459
rect 39806 477461 39866 597211
rect 55998 596733 56058 599390
rect 57102 597141 57162 599390
rect 58206 597413 58266 599390
rect 58203 597412 58269 597413
rect 58203 597348 58204 597412
rect 58268 597348 58269 597412
rect 58203 597347 58269 597348
rect 59494 597141 59554 599390
rect 60598 597277 60658 599390
rect 61702 599390 61828 599450
rect 63128 599450 63188 600100
rect 64216 599450 64276 600100
rect 65440 599450 65500 600100
rect 66528 599450 66588 600100
rect 67616 599450 67676 600100
rect 63128 599390 63234 599450
rect 64216 599390 64338 599450
rect 61702 597549 61762 599390
rect 63174 597549 63234 599390
rect 64278 597549 64338 599390
rect 64646 599390 65500 599450
rect 66486 599390 66588 599450
rect 67590 599390 67676 599450
rect 68296 599450 68356 600100
rect 68704 599450 68764 600100
rect 70064 599450 70124 600100
rect 70744 599450 70804 600100
rect 71288 599450 71348 600100
rect 72376 599450 72436 600100
rect 68296 599390 68386 599450
rect 64646 597549 64706 599390
rect 66486 597549 66546 599390
rect 67590 597549 67650 599390
rect 68326 597549 68386 599390
rect 68694 599390 68764 599450
rect 69982 599390 70124 599450
rect 70718 599390 70804 599450
rect 71270 599390 71348 599450
rect 72374 599390 72436 599450
rect 73464 599450 73524 600100
rect 73600 599450 73660 600100
rect 74552 599450 74612 600100
rect 75912 599450 75972 600100
rect 73464 599390 73538 599450
rect 73600 599390 73722 599450
rect 74552 599390 74642 599450
rect 61699 597548 61765 597549
rect 61699 597484 61700 597548
rect 61764 597484 61765 597548
rect 61699 597483 61765 597484
rect 63171 597548 63237 597549
rect 63171 597484 63172 597548
rect 63236 597484 63237 597548
rect 63171 597483 63237 597484
rect 64275 597548 64341 597549
rect 64275 597484 64276 597548
rect 64340 597484 64341 597548
rect 64275 597483 64341 597484
rect 64643 597548 64709 597549
rect 64643 597484 64644 597548
rect 64708 597484 64709 597548
rect 64643 597483 64709 597484
rect 66483 597548 66549 597549
rect 66483 597484 66484 597548
rect 66548 597484 66549 597548
rect 66483 597483 66549 597484
rect 67587 597548 67653 597549
rect 67587 597484 67588 597548
rect 67652 597484 67653 597548
rect 67587 597483 67653 597484
rect 68323 597548 68389 597549
rect 68323 597484 68324 597548
rect 68388 597484 68389 597548
rect 68323 597483 68389 597484
rect 68694 597413 68754 599390
rect 69982 597549 70042 599390
rect 70718 597549 70778 599390
rect 69979 597548 70045 597549
rect 69979 597484 69980 597548
rect 70044 597484 70045 597548
rect 69979 597483 70045 597484
rect 70715 597548 70781 597549
rect 70715 597484 70716 597548
rect 70780 597484 70781 597548
rect 70715 597483 70781 597484
rect 71270 597413 71330 599390
rect 72374 597413 72434 599390
rect 73478 597549 73538 599390
rect 73662 597549 73722 599390
rect 74582 597549 74642 599390
rect 75870 599390 75972 599450
rect 76048 599450 76108 600100
rect 77000 599450 77060 600100
rect 78088 599450 78148 600100
rect 78496 599450 78556 600100
rect 79448 599450 79508 600100
rect 80672 599450 80732 600100
rect 81080 599450 81140 600100
rect 81760 599450 81820 600100
rect 76048 599390 76114 599450
rect 73475 597548 73541 597549
rect 73475 597484 73476 597548
rect 73540 597484 73541 597548
rect 73475 597483 73541 597484
rect 73659 597548 73725 597549
rect 73659 597484 73660 597548
rect 73724 597484 73725 597548
rect 73659 597483 73725 597484
rect 74579 597548 74645 597549
rect 74579 597484 74580 597548
rect 74644 597484 74645 597548
rect 74579 597483 74645 597484
rect 75870 597413 75930 599390
rect 76054 597549 76114 599390
rect 76974 599390 77060 599450
rect 78078 599390 78148 599450
rect 78446 599390 78556 599450
rect 79366 599390 79508 599450
rect 80654 599390 80732 599450
rect 81022 599390 81140 599450
rect 81758 599390 81820 599450
rect 82848 599450 82908 600100
rect 83528 599450 83588 600100
rect 83936 599450 83996 600100
rect 85296 599450 85356 600100
rect 82848 599390 82922 599450
rect 83528 599390 83658 599450
rect 76051 597548 76117 597549
rect 76051 597484 76052 597548
rect 76116 597484 76117 597548
rect 76051 597483 76117 597484
rect 76974 597413 77034 599390
rect 78078 597549 78138 599390
rect 78446 597549 78506 599390
rect 78075 597548 78141 597549
rect 78075 597484 78076 597548
rect 78140 597484 78141 597548
rect 78075 597483 78141 597484
rect 78443 597548 78509 597549
rect 78443 597484 78444 597548
rect 78508 597484 78509 597548
rect 78443 597483 78509 597484
rect 68691 597412 68757 597413
rect 68691 597348 68692 597412
rect 68756 597348 68757 597412
rect 68691 597347 68757 597348
rect 71267 597412 71333 597413
rect 71267 597348 71268 597412
rect 71332 597348 71333 597412
rect 71267 597347 71333 597348
rect 72371 597412 72437 597413
rect 72371 597348 72372 597412
rect 72436 597348 72437 597412
rect 72371 597347 72437 597348
rect 75867 597412 75933 597413
rect 75867 597348 75868 597412
rect 75932 597348 75933 597412
rect 75867 597347 75933 597348
rect 76971 597412 77037 597413
rect 76971 597348 76972 597412
rect 77036 597348 77037 597412
rect 76971 597347 77037 597348
rect 60595 597276 60661 597277
rect 60595 597212 60596 597276
rect 60660 597212 60661 597276
rect 60595 597211 60661 597212
rect 57099 597140 57165 597141
rect 57099 597076 57100 597140
rect 57164 597076 57165 597140
rect 57099 597075 57165 597076
rect 59491 597140 59557 597141
rect 59491 597076 59492 597140
rect 59556 597076 59557 597140
rect 59491 597075 59557 597076
rect 79366 597005 79426 599390
rect 80654 597005 80714 599390
rect 81022 597549 81082 599390
rect 81019 597548 81085 597549
rect 81019 597484 81020 597548
rect 81084 597484 81085 597548
rect 81019 597483 81085 597484
rect 81758 597277 81818 599390
rect 81755 597276 81821 597277
rect 81755 597212 81756 597276
rect 81820 597212 81821 597276
rect 81755 597211 81821 597212
rect 79363 597004 79429 597005
rect 79363 596940 79364 597004
rect 79428 596940 79429 597004
rect 79363 596939 79429 596940
rect 80651 597004 80717 597005
rect 80651 596940 80652 597004
rect 80716 596940 80717 597004
rect 80651 596939 80717 596940
rect 82862 596869 82922 599390
rect 82859 596868 82925 596869
rect 82859 596804 82860 596868
rect 82924 596804 82925 596868
rect 82859 596803 82925 596804
rect 55995 596732 56061 596733
rect 55995 596668 55996 596732
rect 56060 596668 56061 596732
rect 55995 596667 56061 596668
rect 83598 596461 83658 599390
rect 83782 599390 83996 599450
rect 84334 599390 85356 599450
rect 85976 599450 86036 600100
rect 86384 599450 86444 600100
rect 85976 599390 86050 599450
rect 83782 597413 83842 599390
rect 84334 598770 84394 599390
rect 83966 598710 84394 598770
rect 83966 597549 84026 598710
rect 85990 597549 86050 599390
rect 86358 599390 86444 599450
rect 87608 599450 87668 600100
rect 88288 599450 88348 600100
rect 87608 599390 87706 599450
rect 83963 597548 84029 597549
rect 83963 597484 83964 597548
rect 84028 597484 84029 597548
rect 83963 597483 84029 597484
rect 85987 597548 86053 597549
rect 85987 597484 85988 597548
rect 86052 597484 86053 597548
rect 85987 597483 86053 597484
rect 83779 597412 83845 597413
rect 83779 597348 83780 597412
rect 83844 597348 83845 597412
rect 83779 597347 83845 597348
rect 86358 597277 86418 599390
rect 87646 597277 87706 599390
rect 88198 599390 88348 599450
rect 88696 599450 88756 600100
rect 89784 599450 89844 600100
rect 91008 599450 91068 600100
rect 91144 599450 91204 600100
rect 88696 599390 88810 599450
rect 89784 599390 89914 599450
rect 88198 597549 88258 599390
rect 88195 597548 88261 597549
rect 88195 597484 88196 597548
rect 88260 597484 88261 597548
rect 88195 597483 88261 597484
rect 86355 597276 86421 597277
rect 86355 597212 86356 597276
rect 86420 597212 86421 597276
rect 86355 597211 86421 597212
rect 87643 597276 87709 597277
rect 87643 597212 87644 597276
rect 87708 597212 87709 597276
rect 87643 597211 87709 597212
rect 88750 597141 88810 599390
rect 89854 597141 89914 599390
rect 90958 599390 91068 599450
rect 91142 599390 91204 599450
rect 92232 599450 92292 600100
rect 93320 599450 93380 600100
rect 93592 599450 93652 600100
rect 94408 599586 94468 600100
rect 95768 599586 95828 600100
rect 94408 599526 94514 599586
rect 92232 599390 92306 599450
rect 93320 599390 93410 599450
rect 88747 597140 88813 597141
rect 88747 597076 88748 597140
rect 88812 597076 88813 597140
rect 88747 597075 88813 597076
rect 89851 597140 89917 597141
rect 89851 597076 89852 597140
rect 89916 597076 89917 597140
rect 89851 597075 89917 597076
rect 83595 596460 83661 596461
rect 83595 596396 83596 596460
rect 83660 596396 83661 596460
rect 83595 596395 83661 596396
rect 90958 596325 91018 599390
rect 91142 596461 91202 599390
rect 92246 596597 92306 599390
rect 93350 597549 93410 599390
rect 93534 599390 93652 599450
rect 93534 597549 93594 599390
rect 93347 597548 93413 597549
rect 93347 597484 93348 597548
rect 93412 597484 93413 597548
rect 93347 597483 93413 597484
rect 93531 597548 93597 597549
rect 93531 597484 93532 597548
rect 93596 597484 93597 597548
rect 93531 597483 93597 597484
rect 94454 596597 94514 599526
rect 95742 599526 95828 599586
rect 96040 599586 96100 600100
rect 96992 599586 97052 600100
rect 98080 599586 98140 600100
rect 98488 599586 98548 600100
rect 99168 599586 99228 600100
rect 100936 599586 100996 600100
rect 96040 599526 96170 599586
rect 96992 599526 97090 599586
rect 98080 599526 98194 599586
rect 98488 599526 98562 599586
rect 95742 597277 95802 599526
rect 95739 597276 95805 597277
rect 95739 597212 95740 597276
rect 95804 597212 95805 597276
rect 95739 597211 95805 597212
rect 92243 596596 92309 596597
rect 92243 596532 92244 596596
rect 92308 596532 92309 596596
rect 92243 596531 92309 596532
rect 94451 596596 94517 596597
rect 94451 596532 94452 596596
rect 94516 596532 94517 596596
rect 94451 596531 94517 596532
rect 96110 596461 96170 599526
rect 97030 597141 97090 599526
rect 98134 597413 98194 599526
rect 98131 597412 98197 597413
rect 98131 597348 98132 597412
rect 98196 597348 98197 597412
rect 98131 597347 98197 597348
rect 97027 597140 97093 597141
rect 97027 597076 97028 597140
rect 97092 597076 97093 597140
rect 97027 597075 97093 597076
rect 98502 596461 98562 599526
rect 99054 599526 99228 599586
rect 100894 599526 100996 599586
rect 99054 597277 99114 599526
rect 99051 597276 99117 597277
rect 99051 597212 99052 597276
rect 99116 597212 99117 597276
rect 99051 597211 99117 597212
rect 100894 596733 100954 599526
rect 103520 599450 103580 600100
rect 103286 599390 103580 599450
rect 105968 599450 106028 600100
rect 108280 599450 108340 600100
rect 105968 599390 106106 599450
rect 103286 596869 103346 599390
rect 103283 596868 103349 596869
rect 103283 596804 103284 596868
rect 103348 596804 103349 596868
rect 103283 596803 103349 596804
rect 100891 596732 100957 596733
rect 100891 596668 100892 596732
rect 100956 596668 100957 596732
rect 100891 596667 100957 596668
rect 106046 596597 106106 599390
rect 108254 599390 108340 599450
rect 111000 599450 111060 600100
rect 113448 599450 113508 600100
rect 111000 599390 111074 599450
rect 108254 597413 108314 599390
rect 108251 597412 108317 597413
rect 108251 597348 108252 597412
rect 108316 597348 108317 597412
rect 108251 597347 108317 597348
rect 111014 597005 111074 599390
rect 113406 599390 113508 599450
rect 115896 599450 115956 600100
rect 118480 599450 118540 600100
rect 120928 599450 120988 600100
rect 123512 599450 123572 600100
rect 125960 599450 126020 600100
rect 128544 599450 128604 600100
rect 115896 599390 116042 599450
rect 118480 599390 118618 599450
rect 120928 599390 121010 599450
rect 113406 597277 113466 599390
rect 115982 597413 116042 599390
rect 115979 597412 116045 597413
rect 115979 597348 115980 597412
rect 116044 597348 116045 597412
rect 115979 597347 116045 597348
rect 113403 597276 113469 597277
rect 113403 597212 113404 597276
rect 113468 597212 113469 597276
rect 113403 597211 113469 597212
rect 118558 597005 118618 599390
rect 120950 597413 121010 599390
rect 122606 599390 123572 599450
rect 125918 599390 126020 599450
rect 128494 599390 128604 599450
rect 130992 599450 131052 600100
rect 133440 599450 133500 600100
rect 135888 599450 135948 600100
rect 138472 599450 138532 600100
rect 130992 599390 131130 599450
rect 133440 599390 133522 599450
rect 122606 597549 122666 599390
rect 122603 597548 122669 597549
rect 122603 597484 122604 597548
rect 122668 597484 122669 597548
rect 122603 597483 122669 597484
rect 120947 597412 121013 597413
rect 120947 597348 120948 597412
rect 121012 597348 121013 597412
rect 120947 597347 121013 597348
rect 125918 597141 125978 599390
rect 128494 597549 128554 599390
rect 131070 597549 131130 599390
rect 133462 597549 133522 599390
rect 135854 599390 135948 599450
rect 138430 599390 138532 599450
rect 140920 599450 140980 600100
rect 143368 599450 143428 600100
rect 140920 599390 141066 599450
rect 135854 597549 135914 599390
rect 128491 597548 128557 597549
rect 128491 597484 128492 597548
rect 128556 597484 128557 597548
rect 128491 597483 128557 597484
rect 131067 597548 131133 597549
rect 131067 597484 131068 597548
rect 131132 597484 131133 597548
rect 131067 597483 131133 597484
rect 133459 597548 133525 597549
rect 133459 597484 133460 597548
rect 133524 597484 133525 597548
rect 133459 597483 133525 597484
rect 135851 597548 135917 597549
rect 135851 597484 135852 597548
rect 135916 597484 135917 597548
rect 135851 597483 135917 597484
rect 138430 597141 138490 599390
rect 141006 597549 141066 599390
rect 141926 599390 143428 599450
rect 145952 599450 146012 600100
rect 145952 599390 146034 599450
rect 141003 597548 141069 597549
rect 141003 597484 141004 597548
rect 141068 597484 141069 597548
rect 141003 597483 141069 597484
rect 125915 597140 125981 597141
rect 125915 597076 125916 597140
rect 125980 597076 125981 597140
rect 125915 597075 125981 597076
rect 138427 597140 138493 597141
rect 138427 597076 138428 597140
rect 138492 597076 138493 597140
rect 138427 597075 138493 597076
rect 141926 597005 141986 599390
rect 145974 597549 146034 599390
rect 145971 597548 146037 597549
rect 145971 597484 145972 597548
rect 146036 597484 146037 597548
rect 145971 597483 146037 597484
rect 111011 597004 111077 597005
rect 111011 596940 111012 597004
rect 111076 596940 111077 597004
rect 111011 596939 111077 596940
rect 118555 597004 118621 597005
rect 118555 596940 118556 597004
rect 118620 596940 118621 597004
rect 118555 596939 118621 596940
rect 141923 597004 141989 597005
rect 141923 596940 141924 597004
rect 141988 596940 141989 597004
rect 141923 596939 141989 596940
rect 106043 596596 106109 596597
rect 106043 596532 106044 596596
rect 106108 596532 106109 596596
rect 106043 596531 106109 596532
rect 91139 596460 91205 596461
rect 91139 596396 91140 596460
rect 91204 596396 91205 596460
rect 91139 596395 91205 596396
rect 96107 596460 96173 596461
rect 96107 596396 96108 596460
rect 96172 596396 96173 596460
rect 96107 596395 96173 596396
rect 98499 596460 98565 596461
rect 98499 596396 98500 596460
rect 98564 596396 98565 596460
rect 98499 596395 98565 596396
rect 90955 596324 91021 596325
rect 90955 596260 90956 596324
rect 91020 596260 91021 596324
rect 90955 596259 91021 596260
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 170811 565860 170877 565861
rect 170811 565796 170812 565860
rect 170876 565796 170877 565860
rect 170811 565795 170877 565796
rect 170814 564090 170874 565795
rect 170814 564030 170900 564090
rect 170840 563202 170900 564030
rect 40272 547174 40620 547206
rect 40272 546938 40328 547174
rect 40564 546938 40620 547174
rect 40272 546854 40620 546938
rect 40272 546618 40328 546854
rect 40564 546618 40620 546854
rect 40272 546586 40620 546618
rect 176000 547174 176348 547206
rect 176000 546938 176056 547174
rect 176292 546938 176348 547174
rect 176000 546854 176348 546938
rect 176000 546618 176056 546854
rect 176292 546618 176348 546854
rect 176000 546586 176348 546618
rect 40952 543454 41300 543486
rect 40952 543218 41008 543454
rect 41244 543218 41300 543454
rect 40952 543134 41300 543218
rect 40952 542898 41008 543134
rect 41244 542898 41300 543134
rect 40952 542866 41300 542898
rect 175320 543454 175668 543486
rect 175320 543218 175376 543454
rect 175612 543218 175668 543454
rect 175320 543134 175668 543218
rect 175320 542898 175376 543134
rect 175612 542898 175668 543134
rect 175320 542866 175668 542898
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 40272 511174 40620 511206
rect 40272 510938 40328 511174
rect 40564 510938 40620 511174
rect 40272 510854 40620 510938
rect 40272 510618 40328 510854
rect 40564 510618 40620 510854
rect 40272 510586 40620 510618
rect 176000 511174 176348 511206
rect 176000 510938 176056 511174
rect 176292 510938 176348 511174
rect 176000 510854 176348 510938
rect 176000 510618 176056 510854
rect 176292 510618 176348 510854
rect 176000 510586 176348 510618
rect 40952 507454 41300 507486
rect 40952 507218 41008 507454
rect 41244 507218 41300 507454
rect 40952 507134 41300 507218
rect 40952 506898 41008 507134
rect 41244 506898 41300 507134
rect 40952 506866 41300 506898
rect 175320 507454 175668 507486
rect 175320 507218 175376 507454
rect 175612 507218 175668 507454
rect 175320 507134 175668 507218
rect 175320 506898 175376 507134
rect 175612 506898 175668 507134
rect 175320 506866 175668 506898
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 56056 479637 56116 480080
rect 57144 479770 57204 480080
rect 58232 479770 58292 480080
rect 59592 479770 59652 480080
rect 57102 479710 57204 479770
rect 58206 479710 58292 479770
rect 59494 479710 59652 479770
rect 60544 479770 60604 480080
rect 61768 479770 61828 480080
rect 60544 479710 60658 479770
rect 56053 479636 56119 479637
rect 56053 479572 56054 479636
rect 56118 479572 56119 479636
rect 56053 479571 56119 479572
rect 39803 477460 39869 477461
rect 39803 477396 39804 477460
rect 39868 477396 39869 477460
rect 39803 477395 39869 477396
rect 57102 476781 57162 479710
rect 58206 476917 58266 479710
rect 59494 477325 59554 479710
rect 60598 477461 60658 479710
rect 61702 479710 61828 479770
rect 63128 479770 63188 480080
rect 64216 479770 64276 480080
rect 65440 479770 65500 480080
rect 66528 479770 66588 480080
rect 67616 479770 67676 480080
rect 63128 479710 63234 479770
rect 64216 479710 64338 479770
rect 60595 477460 60661 477461
rect 60595 477396 60596 477460
rect 60660 477396 60661 477460
rect 60595 477395 60661 477396
rect 59491 477324 59557 477325
rect 59491 477260 59492 477324
rect 59556 477260 59557 477324
rect 59491 477259 59557 477260
rect 60598 477053 60658 477395
rect 61702 477325 61762 479710
rect 63174 477461 63234 479710
rect 64278 477461 64338 479710
rect 65382 479710 65500 479770
rect 66486 479710 66588 479770
rect 67590 479710 67676 479770
rect 68296 479770 68356 480080
rect 68704 479770 68764 480080
rect 68296 479710 68386 479770
rect 65382 477461 65442 479710
rect 66486 477461 66546 479710
rect 67590 477461 67650 479710
rect 63171 477460 63237 477461
rect 63171 477396 63172 477460
rect 63236 477396 63237 477460
rect 63171 477395 63237 477396
rect 64275 477460 64341 477461
rect 64275 477396 64276 477460
rect 64340 477396 64341 477460
rect 64275 477395 64341 477396
rect 65379 477460 65445 477461
rect 65379 477396 65380 477460
rect 65444 477396 65445 477460
rect 65379 477395 65445 477396
rect 66483 477460 66549 477461
rect 66483 477396 66484 477460
rect 66548 477396 66549 477460
rect 66483 477395 66549 477396
rect 67587 477460 67653 477461
rect 67587 477396 67588 477460
rect 67652 477396 67653 477460
rect 67587 477395 67653 477396
rect 61699 477324 61765 477325
rect 61699 477260 61700 477324
rect 61764 477260 61765 477324
rect 61699 477259 61765 477260
rect 60595 477052 60661 477053
rect 60595 476988 60596 477052
rect 60660 476988 60661 477052
rect 60595 476987 60661 476988
rect 58203 476916 58269 476917
rect 58203 476852 58204 476916
rect 58268 476852 58269 476916
rect 58203 476851 58269 476852
rect 57099 476780 57165 476781
rect 57099 476716 57100 476780
rect 57164 476716 57165 476780
rect 57099 476715 57165 476716
rect 68326 476237 68386 479710
rect 68694 479710 68764 479770
rect 70064 479770 70124 480080
rect 70744 479770 70804 480080
rect 71288 479770 71348 480080
rect 72376 479770 72436 480080
rect 70064 479710 70226 479770
rect 68694 477461 68754 479710
rect 70166 477461 70226 479710
rect 70718 479710 70804 479770
rect 71270 479710 71348 479770
rect 72374 479710 72436 479770
rect 73464 479770 73524 480080
rect 73600 479770 73660 480080
rect 74552 479770 74612 480080
rect 75912 479770 75972 480080
rect 73464 479710 73538 479770
rect 73600 479710 73722 479770
rect 74552 479710 74642 479770
rect 68691 477460 68757 477461
rect 68691 477396 68692 477460
rect 68756 477396 68757 477460
rect 68691 477395 68757 477396
rect 70163 477460 70229 477461
rect 70163 477396 70164 477460
rect 70228 477396 70229 477460
rect 70163 477395 70229 477396
rect 70718 476237 70778 479710
rect 71270 477461 71330 479710
rect 72374 478685 72434 479710
rect 72371 478684 72437 478685
rect 72371 478620 72372 478684
rect 72436 478620 72437 478684
rect 72371 478619 72437 478620
rect 73478 478549 73538 479710
rect 73475 478548 73541 478549
rect 73475 478484 73476 478548
rect 73540 478484 73541 478548
rect 73475 478483 73541 478484
rect 71267 477460 71333 477461
rect 71267 477396 71268 477460
rect 71332 477396 71333 477460
rect 71267 477395 71333 477396
rect 73662 476237 73722 479710
rect 74582 478685 74642 479710
rect 75870 479710 75972 479770
rect 76048 479770 76108 480080
rect 77000 479770 77060 480080
rect 78088 479770 78148 480080
rect 78496 479770 78556 480080
rect 76048 479710 76114 479770
rect 74579 478684 74645 478685
rect 74579 478620 74580 478684
rect 74644 478620 74645 478684
rect 74579 478619 74645 478620
rect 75870 478413 75930 479710
rect 75867 478412 75933 478413
rect 75867 478348 75868 478412
rect 75932 478348 75933 478412
rect 75867 478347 75933 478348
rect 76054 476237 76114 479710
rect 76974 479710 77060 479770
rect 78078 479710 78148 479770
rect 78446 479710 78556 479770
rect 79448 479770 79508 480080
rect 80672 479770 80732 480080
rect 81080 479770 81140 480080
rect 81760 479770 81820 480080
rect 79448 479710 79610 479770
rect 76974 478549 77034 479710
rect 76971 478548 77037 478549
rect 76971 478484 76972 478548
rect 77036 478484 77037 478548
rect 76971 478483 77037 478484
rect 78078 477461 78138 479710
rect 78075 477460 78141 477461
rect 78075 477396 78076 477460
rect 78140 477396 78141 477460
rect 78075 477395 78141 477396
rect 78446 476237 78506 479710
rect 79550 478277 79610 479710
rect 80654 479710 80732 479770
rect 81022 479710 81140 479770
rect 81758 479710 81820 479770
rect 82848 479770 82908 480080
rect 83528 479770 83588 480080
rect 83936 479770 83996 480080
rect 85296 479770 85356 480080
rect 82848 479710 82922 479770
rect 83528 479710 83658 479770
rect 83936 479710 84026 479770
rect 79547 478276 79613 478277
rect 79547 478212 79548 478276
rect 79612 478212 79613 478276
rect 79547 478211 79613 478212
rect 79550 476373 79610 478211
rect 80654 478141 80714 479710
rect 80651 478140 80717 478141
rect 80651 478076 80652 478140
rect 80716 478076 80717 478140
rect 80651 478075 80717 478076
rect 81022 477461 81082 479710
rect 81758 477461 81818 479710
rect 82862 477461 82922 479710
rect 83598 477461 83658 479710
rect 81019 477460 81085 477461
rect 81019 477396 81020 477460
rect 81084 477396 81085 477460
rect 81019 477395 81085 477396
rect 81755 477460 81821 477461
rect 81755 477396 81756 477460
rect 81820 477396 81821 477460
rect 81755 477395 81821 477396
rect 82859 477460 82925 477461
rect 82859 477396 82860 477460
rect 82924 477396 82925 477460
rect 82859 477395 82925 477396
rect 83595 477460 83661 477461
rect 83595 477396 83596 477460
rect 83660 477396 83661 477460
rect 83595 477395 83661 477396
rect 83966 476645 84026 479710
rect 85254 479710 85356 479770
rect 85976 479770 86036 480080
rect 86384 479770 86444 480080
rect 85976 479710 86050 479770
rect 85254 477461 85314 479710
rect 85990 477461 86050 479710
rect 86358 479710 86444 479770
rect 87608 479770 87668 480080
rect 88288 479770 88348 480080
rect 87608 479710 87706 479770
rect 86358 477597 86418 479710
rect 86355 477596 86421 477597
rect 86355 477532 86356 477596
rect 86420 477532 86421 477596
rect 86355 477531 86421 477532
rect 87646 477461 87706 479710
rect 88198 479710 88348 479770
rect 88696 479770 88756 480080
rect 89784 479770 89844 480080
rect 91008 479770 91068 480080
rect 91144 479770 91204 480080
rect 88696 479710 88810 479770
rect 89784 479710 89914 479770
rect 88198 477461 88258 479710
rect 88750 477461 88810 479710
rect 89854 477461 89914 479710
rect 90958 479710 91068 479770
rect 91142 479710 91204 479770
rect 92232 479770 92292 480080
rect 93320 479770 93380 480080
rect 93592 479770 93652 480080
rect 92232 479710 92306 479770
rect 93320 479710 93410 479770
rect 85251 477460 85317 477461
rect 85251 477396 85252 477460
rect 85316 477396 85317 477460
rect 85251 477395 85317 477396
rect 85987 477460 86053 477461
rect 85987 477396 85988 477460
rect 86052 477396 86053 477460
rect 85987 477395 86053 477396
rect 87643 477460 87709 477461
rect 87643 477396 87644 477460
rect 87708 477396 87709 477460
rect 87643 477395 87709 477396
rect 88195 477460 88261 477461
rect 88195 477396 88196 477460
rect 88260 477396 88261 477460
rect 88195 477395 88261 477396
rect 88747 477460 88813 477461
rect 88747 477396 88748 477460
rect 88812 477396 88813 477460
rect 88747 477395 88813 477396
rect 89851 477460 89917 477461
rect 89851 477396 89852 477460
rect 89916 477396 89917 477460
rect 89851 477395 89917 477396
rect 83963 476644 84029 476645
rect 83963 476580 83964 476644
rect 84028 476580 84029 476644
rect 83963 476579 84029 476580
rect 90958 476509 91018 479710
rect 91142 477461 91202 479710
rect 92246 477461 92306 479710
rect 93350 477461 93410 479710
rect 93534 479710 93652 479770
rect 94408 479770 94468 480080
rect 95768 479770 95828 480080
rect 94408 479710 94514 479770
rect 91139 477460 91205 477461
rect 91139 477396 91140 477460
rect 91204 477396 91205 477460
rect 91139 477395 91205 477396
rect 92243 477460 92309 477461
rect 92243 477396 92244 477460
rect 92308 477396 92309 477460
rect 92243 477395 92309 477396
rect 93347 477460 93413 477461
rect 93347 477396 93348 477460
rect 93412 477396 93413 477460
rect 93347 477395 93413 477396
rect 93534 476509 93594 479710
rect 94454 477461 94514 479710
rect 95742 479710 95828 479770
rect 96040 479770 96100 480080
rect 96992 479770 97052 480080
rect 98080 479770 98140 480080
rect 98488 479770 98548 480080
rect 99168 479770 99228 480080
rect 100936 479770 100996 480080
rect 103520 479770 103580 480080
rect 96040 479710 96170 479770
rect 96992 479710 97090 479770
rect 98080 479710 98194 479770
rect 98488 479710 98562 479770
rect 95742 477461 95802 479710
rect 94451 477460 94517 477461
rect 94451 477396 94452 477460
rect 94516 477396 94517 477460
rect 94451 477395 94517 477396
rect 95739 477460 95805 477461
rect 95739 477396 95740 477460
rect 95804 477396 95805 477460
rect 95739 477395 95805 477396
rect 90955 476508 91021 476509
rect 90955 476444 90956 476508
rect 91020 476444 91021 476508
rect 90955 476443 91021 476444
rect 93531 476508 93597 476509
rect 93531 476444 93532 476508
rect 93596 476444 93597 476508
rect 93531 476443 93597 476444
rect 79547 476372 79613 476373
rect 79547 476308 79548 476372
rect 79612 476308 79613 476372
rect 79547 476307 79613 476308
rect 96110 476237 96170 479710
rect 97030 477461 97090 479710
rect 97027 477460 97093 477461
rect 97027 477396 97028 477460
rect 97092 477396 97093 477460
rect 97027 477395 97093 477396
rect 98134 476373 98194 479710
rect 98131 476372 98197 476373
rect 98131 476308 98132 476372
rect 98196 476308 98197 476372
rect 98131 476307 98197 476308
rect 98502 476237 98562 479710
rect 99054 479710 99228 479770
rect 100894 479710 100996 479770
rect 103286 479710 103580 479770
rect 105968 479770 106028 480080
rect 108280 479770 108340 480080
rect 105968 479710 106106 479770
rect 99054 477461 99114 479710
rect 99051 477460 99117 477461
rect 99051 477396 99052 477460
rect 99116 477396 99117 477460
rect 99051 477395 99117 477396
rect 99054 476509 99114 477395
rect 99051 476508 99117 476509
rect 99051 476444 99052 476508
rect 99116 476444 99117 476508
rect 99051 476443 99117 476444
rect 100894 476237 100954 479710
rect 103286 476642 103346 479710
rect 103286 476582 103714 476642
rect 103654 476237 103714 476582
rect 106046 476237 106106 479710
rect 108254 479710 108340 479770
rect 111000 479770 111060 480080
rect 113448 479770 113508 480080
rect 111000 479710 111074 479770
rect 108254 476237 108314 479710
rect 111014 476237 111074 479710
rect 113406 479710 113508 479770
rect 115896 479770 115956 480080
rect 118480 479770 118540 480080
rect 120928 479770 120988 480080
rect 123512 479770 123572 480080
rect 125960 479770 126020 480080
rect 128544 479770 128604 480080
rect 115896 479710 116042 479770
rect 118480 479710 118618 479770
rect 120928 479710 121010 479770
rect 123512 479710 123586 479770
rect 113406 476237 113466 479710
rect 115982 476237 116042 479710
rect 118558 476237 118618 479710
rect 120950 476237 121010 479710
rect 123526 476237 123586 479710
rect 125918 479710 126020 479770
rect 128494 479710 128604 479770
rect 130992 479770 131052 480080
rect 133440 479770 133500 480080
rect 135888 479770 135948 480080
rect 138472 479770 138532 480080
rect 130992 479710 131130 479770
rect 133440 479710 133522 479770
rect 125918 476237 125978 479710
rect 128494 476237 128554 479710
rect 131070 476237 131130 479710
rect 133462 476237 133522 479710
rect 135854 479710 135948 479770
rect 138430 479710 138532 479770
rect 140920 479770 140980 480080
rect 143368 479770 143428 480080
rect 145952 479770 146012 480080
rect 140920 479710 141066 479770
rect 143368 479710 143458 479770
rect 145952 479710 146034 479770
rect 135854 476237 135914 479710
rect 138430 476237 138490 479710
rect 141006 476237 141066 479710
rect 143398 476237 143458 479710
rect 145974 476237 146034 479710
rect 68323 476236 68389 476237
rect 68323 476172 68324 476236
rect 68388 476172 68389 476236
rect 68323 476171 68389 476172
rect 70715 476236 70781 476237
rect 70715 476172 70716 476236
rect 70780 476172 70781 476236
rect 70715 476171 70781 476172
rect 73659 476236 73725 476237
rect 73659 476172 73660 476236
rect 73724 476172 73725 476236
rect 73659 476171 73725 476172
rect 76051 476236 76117 476237
rect 76051 476172 76052 476236
rect 76116 476172 76117 476236
rect 76051 476171 76117 476172
rect 78443 476236 78509 476237
rect 78443 476172 78444 476236
rect 78508 476172 78509 476236
rect 78443 476171 78509 476172
rect 96107 476236 96173 476237
rect 96107 476172 96108 476236
rect 96172 476172 96173 476236
rect 96107 476171 96173 476172
rect 98499 476236 98565 476237
rect 98499 476172 98500 476236
rect 98564 476172 98565 476236
rect 98499 476171 98565 476172
rect 100891 476236 100957 476237
rect 100891 476172 100892 476236
rect 100956 476172 100957 476236
rect 100891 476171 100957 476172
rect 103651 476236 103717 476237
rect 103651 476172 103652 476236
rect 103716 476172 103717 476236
rect 103651 476171 103717 476172
rect 106043 476236 106109 476237
rect 106043 476172 106044 476236
rect 106108 476172 106109 476236
rect 106043 476171 106109 476172
rect 108251 476236 108317 476237
rect 108251 476172 108252 476236
rect 108316 476172 108317 476236
rect 108251 476171 108317 476172
rect 111011 476236 111077 476237
rect 111011 476172 111012 476236
rect 111076 476172 111077 476236
rect 111011 476171 111077 476172
rect 113403 476236 113469 476237
rect 113403 476172 113404 476236
rect 113468 476172 113469 476236
rect 113403 476171 113469 476172
rect 115979 476236 116045 476237
rect 115979 476172 115980 476236
rect 116044 476172 116045 476236
rect 115979 476171 116045 476172
rect 118555 476236 118621 476237
rect 118555 476172 118556 476236
rect 118620 476172 118621 476236
rect 118555 476171 118621 476172
rect 120947 476236 121013 476237
rect 120947 476172 120948 476236
rect 121012 476172 121013 476236
rect 120947 476171 121013 476172
rect 123523 476236 123589 476237
rect 123523 476172 123524 476236
rect 123588 476172 123589 476236
rect 123523 476171 123589 476172
rect 125915 476236 125981 476237
rect 125915 476172 125916 476236
rect 125980 476172 125981 476236
rect 125915 476171 125981 476172
rect 128491 476236 128557 476237
rect 128491 476172 128492 476236
rect 128556 476172 128557 476236
rect 128491 476171 128557 476172
rect 131067 476236 131133 476237
rect 131067 476172 131068 476236
rect 131132 476172 131133 476236
rect 131067 476171 131133 476172
rect 133459 476236 133525 476237
rect 133459 476172 133460 476236
rect 133524 476172 133525 476236
rect 133459 476171 133525 476172
rect 135851 476236 135917 476237
rect 135851 476172 135852 476236
rect 135916 476172 135917 476236
rect 135851 476171 135917 476172
rect 138427 476236 138493 476237
rect 138427 476172 138428 476236
rect 138492 476172 138493 476236
rect 138427 476171 138493 476172
rect 141003 476236 141069 476237
rect 141003 476172 141004 476236
rect 141068 476172 141069 476236
rect 141003 476171 141069 476172
rect 143395 476236 143461 476237
rect 143395 476172 143396 476236
rect 143460 476172 143461 476236
rect 143395 476171 143461 476172
rect 145971 476236 146037 476237
rect 145971 476172 145972 476236
rect 146036 476172 146037 476236
rect 145971 476171 146037 476172
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 170811 445772 170877 445773
rect 170811 445708 170812 445772
rect 170876 445708 170877 445772
rect 170811 445707 170877 445708
rect 170814 443730 170874 445707
rect 170814 443670 170900 443730
rect 170840 443202 170900 443670
rect 40272 439174 40620 439206
rect 40272 438938 40328 439174
rect 40564 438938 40620 439174
rect 40272 438854 40620 438938
rect 40272 438618 40328 438854
rect 40564 438618 40620 438854
rect 40272 438586 40620 438618
rect 176000 439174 176348 439206
rect 176000 438938 176056 439174
rect 176292 438938 176348 439174
rect 176000 438854 176348 438938
rect 176000 438618 176056 438854
rect 176292 438618 176348 438854
rect 176000 438586 176348 438618
rect 40952 435454 41300 435486
rect 40952 435218 41008 435454
rect 41244 435218 41300 435454
rect 40952 435134 41300 435218
rect 40952 434898 41008 435134
rect 41244 434898 41300 435134
rect 40952 434866 41300 434898
rect 175320 435454 175668 435486
rect 175320 435218 175376 435454
rect 175612 435218 175668 435454
rect 175320 435134 175668 435218
rect 175320 434898 175376 435134
rect 175612 434898 175668 435134
rect 175320 434866 175668 434898
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 40272 403174 40620 403206
rect 40272 402938 40328 403174
rect 40564 402938 40620 403174
rect 40272 402854 40620 402938
rect 40272 402618 40328 402854
rect 40564 402618 40620 402854
rect 40272 402586 40620 402618
rect 176000 403174 176348 403206
rect 176000 402938 176056 403174
rect 176292 402938 176348 403174
rect 176000 402854 176348 402938
rect 176000 402618 176056 402854
rect 176292 402618 176348 402854
rect 176000 402586 176348 402618
rect 40952 399454 41300 399486
rect 40952 399218 41008 399454
rect 41244 399218 41300 399454
rect 40952 399134 41300 399218
rect 40952 398898 41008 399134
rect 41244 398898 41300 399134
rect 40952 398866 41300 398898
rect 175320 399454 175668 399486
rect 175320 399218 175376 399454
rect 175612 399218 175668 399454
rect 175320 399134 175668 399218
rect 175320 398898 175376 399134
rect 175612 398898 175668 399134
rect 175320 398866 175668 398898
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 40272 367174 40620 367206
rect 40272 366938 40328 367174
rect 40564 366938 40620 367174
rect 40272 366854 40620 366938
rect 40272 366618 40328 366854
rect 40564 366618 40620 366854
rect 40272 366586 40620 366618
rect 176000 367174 176348 367206
rect 176000 366938 176056 367174
rect 176292 366938 176348 367174
rect 176000 366854 176348 366938
rect 176000 366618 176056 366854
rect 176292 366618 176348 366854
rect 176000 366586 176348 366618
rect 40952 363454 41300 363486
rect 40952 363218 41008 363454
rect 41244 363218 41300 363454
rect 40952 363134 41300 363218
rect 40952 362898 41008 363134
rect 41244 362898 41300 363134
rect 40952 362866 41300 362898
rect 175320 363454 175668 363486
rect 175320 363218 175376 363454
rect 175612 363218 175668 363454
rect 175320 363134 175668 363218
rect 175320 362898 175376 363134
rect 175612 362898 175668 363134
rect 175320 362866 175668 362898
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 56056 359410 56116 360060
rect 57144 359410 57204 360060
rect 58232 359410 58292 360060
rect 55998 359350 56116 359410
rect 57102 359350 57204 359410
rect 58206 359350 58292 359410
rect 59592 359410 59652 360060
rect 60544 359410 60604 360060
rect 61768 359410 61828 360060
rect 63128 359410 63188 360060
rect 64216 359410 64276 360060
rect 65440 359410 65500 360060
rect 66528 359410 66588 360060
rect 67616 359410 67676 360060
rect 59592 359350 59738 359410
rect 60544 359350 60658 359410
rect 61768 359350 61946 359410
rect 63128 359350 63234 359410
rect 64216 359350 64338 359410
rect 41514 331174 42134 358064
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 38883 304196 38949 304197
rect 38883 304132 38884 304196
rect 38948 304132 38949 304196
rect 38883 304131 38949 304132
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 334894 45854 358064
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 338614 49574 358064
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 342334 53294 358064
rect 55998 357373 56058 359350
rect 55995 357372 56061 357373
rect 55995 357308 55996 357372
rect 56060 357308 56061 357372
rect 55995 357307 56061 357308
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 126334 53294 161778
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52674 90334 53294 125778
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52674 54334 53294 89778
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 346054 57014 358064
rect 57102 357237 57162 359350
rect 58206 357373 58266 359350
rect 59678 357373 59738 359350
rect 60598 358189 60658 359350
rect 60595 358188 60661 358189
rect 60595 358124 60596 358188
rect 60660 358124 60661 358188
rect 60595 358123 60661 358124
rect 58203 357372 58269 357373
rect 58203 357308 58204 357372
rect 58268 357308 58269 357372
rect 58203 357307 58269 357308
rect 59675 357372 59741 357373
rect 59675 357308 59676 357372
rect 59740 357308 59741 357372
rect 59675 357307 59741 357308
rect 57099 357236 57165 357237
rect 57099 357172 57100 357236
rect 57164 357172 57165 357236
rect 57099 357171 57165 357172
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 56394 274054 57014 309498
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 56394 238054 57014 273498
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 56394 130054 57014 165498
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 56394 94054 57014 129498
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 56394 58054 57014 93498
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 349774 60734 357940
rect 61886 357373 61946 359350
rect 63174 357373 63234 359350
rect 64278 358189 64338 359350
rect 64646 359350 65500 359410
rect 66486 359350 66588 359410
rect 67590 359350 67676 359410
rect 68296 359410 68356 360060
rect 68704 359410 68764 360060
rect 68296 359350 68386 359410
rect 64275 358188 64341 358189
rect 64275 358124 64276 358188
rect 64340 358124 64341 358188
rect 64275 358123 64341 358124
rect 61883 357372 61949 357373
rect 61883 357308 61884 357372
rect 61948 357308 61949 357372
rect 61883 357307 61949 357308
rect 63171 357372 63237 357373
rect 63171 357308 63172 357372
rect 63236 357308 63237 357372
rect 63171 357307 63237 357308
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 277774 60734 313218
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 241774 60734 277218
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 60114 205774 60734 241218
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 60114 169774 60734 205218
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 60114 133774 60734 169218
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 60114 97774 60734 133218
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 60114 61774 60734 97218
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 60114 25774 60734 61218
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 353494 64454 357940
rect 64646 356149 64706 359350
rect 66486 357373 66546 359350
rect 66483 357372 66549 357373
rect 66483 357308 66484 357372
rect 66548 357308 66549 357372
rect 66483 357307 66549 357308
rect 67590 356149 67650 359350
rect 68326 357101 68386 359350
rect 68694 359350 68764 359410
rect 70064 359410 70124 360060
rect 70744 359410 70804 360060
rect 71288 359410 71348 360060
rect 72376 359410 72436 360060
rect 73464 359410 73524 360060
rect 70064 359350 70226 359410
rect 68694 357373 68754 359350
rect 70166 357373 70226 359350
rect 70718 359350 70804 359410
rect 71270 359350 71348 359410
rect 72374 359350 72436 359410
rect 73294 359350 73524 359410
rect 73600 359410 73660 360060
rect 74552 359410 74612 360060
rect 75912 359410 75972 360060
rect 73600 359350 73722 359410
rect 74552 359350 74642 359410
rect 68691 357372 68757 357373
rect 68691 357308 68692 357372
rect 68756 357308 68757 357372
rect 68691 357307 68757 357308
rect 70163 357372 70229 357373
rect 70163 357308 70164 357372
rect 70228 357308 70229 357372
rect 70163 357307 70229 357308
rect 70718 357237 70778 359350
rect 71270 357373 71330 359350
rect 72374 357373 72434 359350
rect 71267 357372 71333 357373
rect 71267 357308 71268 357372
rect 71332 357308 71333 357372
rect 71267 357307 71333 357308
rect 72371 357372 72437 357373
rect 72371 357308 72372 357372
rect 72436 357308 72437 357372
rect 72371 357307 72437 357308
rect 73294 357237 73354 359350
rect 73662 358730 73722 359350
rect 73478 358670 73722 358730
rect 73478 357373 73538 358670
rect 73475 357372 73541 357373
rect 73475 357308 73476 357372
rect 73540 357308 73541 357372
rect 73475 357307 73541 357308
rect 70715 357236 70781 357237
rect 70715 357172 70716 357236
rect 70780 357172 70781 357236
rect 70715 357171 70781 357172
rect 73291 357236 73357 357237
rect 73291 357172 73292 357236
rect 73356 357172 73357 357236
rect 73291 357171 73357 357172
rect 68323 357100 68389 357101
rect 68323 357036 68324 357100
rect 68388 357036 68389 357100
rect 68323 357035 68389 357036
rect 64643 356148 64709 356149
rect 64643 356084 64644 356148
rect 64708 356084 64709 356148
rect 64643 356083 64709 356084
rect 67587 356148 67653 356149
rect 67587 356084 67588 356148
rect 67652 356084 67653 356148
rect 67587 356083 67653 356084
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 317494 64454 352938
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 63834 281494 64454 316938
rect 63834 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 64454 281494
rect 63834 281174 64454 281258
rect 63834 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 64454 281174
rect 63834 245494 64454 280938
rect 63834 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 64454 245494
rect 63834 245174 64454 245258
rect 63834 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 64454 245174
rect 63834 209494 64454 244938
rect 63834 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 64454 209494
rect 63834 209174 64454 209258
rect 63834 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 64454 209174
rect 63834 173494 64454 208938
rect 63834 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 64454 173494
rect 63834 173174 64454 173258
rect 63834 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 64454 173174
rect 63834 137494 64454 172938
rect 63834 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 64454 137494
rect 63834 137174 64454 137258
rect 63834 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 64454 137174
rect 63834 101494 64454 136938
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 63834 65494 64454 100938
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 63834 29494 64454 64938
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 327454 74414 358064
rect 74582 357373 74642 359350
rect 75870 359350 75972 359410
rect 76048 359410 76108 360060
rect 77000 359410 77060 360060
rect 76048 359350 76114 359410
rect 74579 357372 74645 357373
rect 74579 357308 74580 357372
rect 74644 357308 74645 357372
rect 74579 357307 74645 357308
rect 75870 357237 75930 359350
rect 75867 357236 75933 357237
rect 75867 357172 75868 357236
rect 75932 357172 75933 357236
rect 75867 357171 75933 357172
rect 76054 356421 76114 359350
rect 76974 359350 77060 359410
rect 78088 359410 78148 360060
rect 78496 359410 78556 360060
rect 78088 359350 78322 359410
rect 76974 357373 77034 359350
rect 76971 357372 77037 357373
rect 76971 357308 76972 357372
rect 77036 357308 77037 357372
rect 76971 357307 77037 357308
rect 76051 356420 76117 356421
rect 76051 356356 76052 356420
rect 76116 356356 76117 356420
rect 76051 356355 76117 356356
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 331174 78134 357940
rect 78262 357237 78322 359350
rect 78446 359350 78556 359410
rect 79448 359410 79508 360060
rect 80672 359410 80732 360060
rect 81080 359410 81140 360060
rect 79448 359350 79610 359410
rect 78446 357373 78506 359350
rect 79550 357373 79610 359350
rect 80654 359350 80732 359410
rect 81022 359350 81140 359410
rect 83528 359410 83588 360060
rect 85976 359410 86036 360060
rect 88288 359410 88348 360060
rect 91008 359410 91068 360060
rect 93592 359410 93652 360060
rect 96040 359410 96100 360060
rect 83528 359350 83658 359410
rect 85976 359350 86050 359410
rect 78443 357372 78509 357373
rect 78443 357308 78444 357372
rect 78508 357308 78509 357372
rect 78443 357307 78509 357308
rect 79547 357372 79613 357373
rect 79547 357308 79548 357372
rect 79612 357308 79613 357372
rect 79547 357307 79613 357308
rect 80654 357237 80714 359350
rect 81022 357373 81082 359350
rect 81019 357372 81085 357373
rect 81019 357308 81020 357372
rect 81084 357308 81085 357372
rect 81019 357307 81085 357308
rect 78259 357236 78325 357237
rect 78259 357172 78260 357236
rect 78324 357172 78325 357236
rect 78259 357171 78325 357172
rect 80651 357236 80717 357237
rect 80651 357172 80652 357236
rect 80716 357172 80717 357236
rect 80651 357171 80717 357172
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 334894 81854 357940
rect 83598 356693 83658 359350
rect 83595 356692 83661 356693
rect 83595 356628 83596 356692
rect 83660 356628 83661 356692
rect 83595 356627 83661 356628
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 338614 85574 357940
rect 85990 357373 86050 359350
rect 88198 359350 88348 359410
rect 90958 359350 91068 359410
rect 93534 359350 93652 359410
rect 95926 359350 96100 359410
rect 98488 359410 98548 360060
rect 100936 359410 100996 360060
rect 103520 359410 103580 360060
rect 98488 359350 98562 359410
rect 88198 357373 88258 359350
rect 85987 357372 86053 357373
rect 85987 357308 85988 357372
rect 86052 357308 86053 357372
rect 85987 357307 86053 357308
rect 88195 357372 88261 357373
rect 88195 357308 88196 357372
rect 88260 357308 88261 357372
rect 88195 357307 88261 357308
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 342334 89294 357940
rect 90958 357373 91018 359350
rect 90955 357372 91021 357373
rect 90955 357308 90956 357372
rect 91020 357308 91021 357372
rect 90955 357307 91021 357308
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 306334 89294 341778
rect 88674 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 89294 306334
rect 88674 306014 89294 306098
rect 88674 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 89294 306014
rect 88674 270334 89294 305778
rect 88674 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 89294 270334
rect 88674 270014 89294 270098
rect 88674 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 89294 270014
rect 88674 234334 89294 269778
rect 88674 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 89294 234334
rect 88674 234014 89294 234098
rect 88674 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 89294 234014
rect 88674 198334 89294 233778
rect 88674 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 89294 198334
rect 88674 198014 89294 198098
rect 88674 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 89294 198014
rect 88674 162334 89294 197778
rect 88674 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 89294 162334
rect 88674 162014 89294 162098
rect 88674 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 89294 162014
rect 88674 126334 89294 161778
rect 88674 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 89294 126334
rect 88674 126014 89294 126098
rect 88674 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 89294 126014
rect 88674 90334 89294 125778
rect 88674 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 89294 90334
rect 88674 90014 89294 90098
rect 88674 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 89294 90014
rect 88674 54334 89294 89778
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 346054 93014 358064
rect 93534 357373 93594 359350
rect 95926 357373 95986 359350
rect 93531 357372 93597 357373
rect 93531 357308 93532 357372
rect 93596 357308 93597 357372
rect 93531 357307 93597 357308
rect 95923 357372 95989 357373
rect 95923 357308 95924 357372
rect 95988 357308 95989 357372
rect 95923 357307 95989 357308
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 310054 93014 345498
rect 92394 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 93014 310054
rect 92394 309734 93014 309818
rect 92394 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 93014 309734
rect 92394 274054 93014 309498
rect 92394 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 93014 274054
rect 92394 273734 93014 273818
rect 92394 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 93014 273734
rect 92394 238054 93014 273498
rect 92394 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 93014 238054
rect 92394 237734 93014 237818
rect 92394 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 93014 237734
rect 92394 202054 93014 237498
rect 92394 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 93014 202054
rect 92394 201734 93014 201818
rect 92394 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 93014 201734
rect 92394 166054 93014 201498
rect 92394 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 93014 166054
rect 92394 165734 93014 165818
rect 92394 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 93014 165734
rect 92394 130054 93014 165498
rect 92394 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 93014 130054
rect 92394 129734 93014 129818
rect 92394 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 93014 129734
rect 92394 94054 93014 129498
rect 92394 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 93014 94054
rect 92394 93734 93014 93818
rect 92394 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 93014 93734
rect 92394 58054 93014 93498
rect 92394 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 93014 58054
rect 92394 57734 93014 57818
rect 92394 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 93014 57734
rect 92394 22054 93014 57498
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 349774 96734 357940
rect 98502 357373 98562 359350
rect 100894 359350 100996 359410
rect 103286 359350 103580 359410
rect 105968 359410 106028 360060
rect 105968 359350 106106 359410
rect 98499 357372 98565 357373
rect 98499 357308 98500 357372
rect 98564 357308 98565 357372
rect 98499 357307 98565 357308
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 313774 96734 349218
rect 96114 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 96734 313774
rect 96114 313454 96734 313538
rect 96114 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 96734 313454
rect 96114 277774 96734 313218
rect 96114 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 96734 277774
rect 96114 277454 96734 277538
rect 96114 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 96734 277454
rect 96114 241774 96734 277218
rect 96114 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 96734 241774
rect 96114 241454 96734 241538
rect 96114 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 96734 241454
rect 96114 205774 96734 241218
rect 96114 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 96734 205774
rect 96114 205454 96734 205538
rect 96114 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 96734 205454
rect 96114 169774 96734 205218
rect 96114 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 96734 169774
rect 96114 169454 96734 169538
rect 96114 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 96734 169454
rect 96114 133774 96734 169218
rect 96114 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 96734 133774
rect 96114 133454 96734 133538
rect 96114 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 96734 133454
rect 96114 97774 96734 133218
rect 96114 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 96734 97774
rect 96114 97454 96734 97538
rect 96114 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 96734 97454
rect 96114 61774 96734 97218
rect 96114 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 96734 61774
rect 96114 61454 96734 61538
rect 96114 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 96734 61454
rect 96114 25774 96734 61218
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 353494 100454 358064
rect 100894 357373 100954 359350
rect 100891 357372 100957 357373
rect 100891 357308 100892 357372
rect 100956 357308 100957 357372
rect 100891 357307 100957 357308
rect 103286 356149 103346 359350
rect 106046 357373 106106 359350
rect 106043 357372 106109 357373
rect 106043 357308 106044 357372
rect 106108 357308 106109 357372
rect 106043 357307 106109 357308
rect 103283 356148 103349 356149
rect 103283 356084 103284 356148
rect 103348 356084 103349 356148
rect 103283 356083 103349 356084
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 317494 100454 352938
rect 99834 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 100454 317494
rect 99834 317174 100454 317258
rect 99834 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 100454 317174
rect 99834 281494 100454 316938
rect 99834 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 100454 281494
rect 99834 281174 100454 281258
rect 99834 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 100454 281174
rect 99834 245494 100454 280938
rect 99834 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 100454 245494
rect 99834 245174 100454 245258
rect 99834 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 100454 245174
rect 99834 209494 100454 244938
rect 99834 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 100454 209494
rect 99834 209174 100454 209258
rect 99834 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 100454 209174
rect 99834 173494 100454 208938
rect 99834 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 100454 173494
rect 99834 173174 100454 173258
rect 99834 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 100454 173174
rect 99834 137494 100454 172938
rect 99834 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 100454 137494
rect 99834 137174 100454 137258
rect 99834 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 100454 137174
rect 99834 101494 100454 136938
rect 99834 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 100454 101494
rect 99834 101174 100454 101258
rect 99834 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 100454 101174
rect 99834 65494 100454 100938
rect 99834 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 100454 65494
rect 99834 65174 100454 65258
rect 99834 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 100454 65174
rect 99834 29494 100454 64938
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 327454 110414 358064
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 331174 114134 357940
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 334894 117854 358064
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 338614 121574 357940
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 124674 342334 125294 358064
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 123707 279580 123773 279581
rect 123707 279516 123708 279580
rect 123772 279516 123773 279580
rect 123707 279515 123773 279516
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 123710 31789 123770 279515
rect 123891 279308 123957 279309
rect 123891 279244 123892 279308
rect 123956 279244 123957 279308
rect 123891 279243 123957 279244
rect 123707 31788 123773 31789
rect 123707 31724 123708 31788
rect 123772 31724 123773 31788
rect 123707 31723 123773 31724
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 123894 7581 123954 279243
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 124208 183454 124528 183486
rect 124208 183218 124250 183454
rect 124486 183218 124528 183454
rect 124208 183134 124528 183218
rect 124208 182898 124250 183134
rect 124486 182898 124528 183134
rect 124208 182866 124528 182898
rect 124674 162334 125294 197778
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 124208 147454 124528 147486
rect 124208 147218 124250 147454
rect 124486 147218 124528 147454
rect 124208 147134 124528 147218
rect 124208 146898 124250 147134
rect 124486 146898 124528 147134
rect 124208 146866 124528 146898
rect 124674 126334 125294 161778
rect 124674 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 125294 126334
rect 124674 126014 125294 126098
rect 124674 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 125294 126014
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 124674 90334 125294 125778
rect 124674 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 125294 90334
rect 124674 90014 125294 90098
rect 124674 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 125294 90014
rect 124674 54334 125294 89778
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 123891 7580 123957 7581
rect 123891 7516 123892 7580
rect 123956 7516 123957 7580
rect 123891 7515 123957 7516
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 346054 129014 357940
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 166054 129014 201498
rect 128394 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 129014 166054
rect 128394 165734 129014 165818
rect 128394 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 129014 165734
rect 128394 130054 129014 165498
rect 128394 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 129014 130054
rect 128394 129734 129014 129818
rect 128394 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 129014 129734
rect 128394 94054 129014 129498
rect 128394 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 129014 94054
rect 128394 93734 129014 93818
rect 128394 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 129014 93734
rect 128394 58054 129014 93498
rect 128394 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 129014 58054
rect 128394 57734 129014 57818
rect 128394 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 129014 57734
rect 128394 22054 129014 57498
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 349774 132734 358064
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 169774 132734 205218
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 132114 169454 132734 169538
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 132114 133774 132734 169218
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 132114 97774 132734 133218
rect 132114 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 132734 97774
rect 132114 97454 132734 97538
rect 132114 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 132734 97454
rect 132114 61774 132734 97218
rect 132114 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 132734 61774
rect 132114 61454 132734 61538
rect 132114 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 132734 61454
rect 132114 25774 132734 61218
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 353494 136454 357940
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 145794 327454 146414 357940
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 139568 259174 139888 259206
rect 139568 258938 139610 259174
rect 139846 258938 139888 259174
rect 139568 258854 139888 258938
rect 139568 258618 139610 258854
rect 139846 258618 139888 258854
rect 139568 258586 139888 258618
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 139568 223174 139888 223206
rect 139568 222938 139610 223174
rect 139846 222938 139888 223174
rect 139568 222854 139888 222938
rect 139568 222618 139610 222854
rect 139846 222618 139888 222854
rect 139568 222586 139888 222618
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 135834 173494 136454 208938
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 139568 187174 139888 187206
rect 139568 186938 139610 187174
rect 139846 186938 139888 187174
rect 139568 186854 139888 186938
rect 139568 186618 139610 186854
rect 139846 186618 139888 186854
rect 139568 186586 139888 186618
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 135834 137494 136454 172938
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 139568 151174 139888 151206
rect 139568 150938 139610 151174
rect 139846 150938 139888 151174
rect 139568 150854 139888 150938
rect 139568 150618 139610 150854
rect 139846 150618 139888 150854
rect 139568 150586 139888 150618
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 135834 101494 136454 136938
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 139568 115174 139888 115206
rect 139568 114938 139610 115174
rect 139846 114938 139888 115174
rect 139568 114854 139888 114938
rect 139568 114618 139610 114854
rect 139846 114618 139888 114854
rect 139568 114586 139888 114618
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 135834 65494 136454 100938
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 135834 29494 136454 64938
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 331174 150134 358064
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 334894 153854 358064
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 156954 338614 157574 358064
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 154928 183454 155248 183486
rect 154928 183218 154970 183454
rect 155206 183218 155248 183454
rect 154928 183134 155248 183218
rect 154928 182898 154970 183134
rect 155206 182898 155248 183134
rect 154928 182866 155248 182898
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 154928 147454 155248 147486
rect 154928 147218 154970 147454
rect 155206 147218 155248 147454
rect 154928 147134 155248 147218
rect 154928 146898 154970 147134
rect 155206 146898 155248 147134
rect 154928 146866 155248 146898
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 342334 161294 358064
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 160674 270334 161294 305778
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 346054 165014 358064
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 349774 168734 358064
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 168114 241774 168734 277218
rect 171834 353494 172454 358064
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 170288 259174 170608 259206
rect 170288 258938 170330 259174
rect 170566 258938 170608 259174
rect 170288 258854 170608 258938
rect 170288 258618 170330 258854
rect 170566 258618 170608 258854
rect 170288 258586 170608 258618
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 171834 245494 172454 280938
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 170288 223174 170608 223206
rect 170288 222938 170330 223174
rect 170566 222938 170608 223174
rect 170288 222854 170608 222938
rect 170288 222618 170330 222854
rect 170566 222618 170608 222854
rect 170288 222586 170608 222618
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 170288 187174 170608 187206
rect 170288 186938 170330 187174
rect 170566 186938 170608 187174
rect 170288 186854 170608 186938
rect 170288 186618 170330 186854
rect 170566 186618 170608 186854
rect 170288 186586 170608 186618
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 170288 151174 170608 151206
rect 170288 150938 170330 151174
rect 170566 150938 170608 151174
rect 170288 150854 170608 150938
rect 170288 150618 170330 150854
rect 170566 150618 170608 150854
rect 170288 150586 170608 150618
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 170288 115174 170608 115206
rect 170288 114938 170330 115174
rect 170566 114938 170608 115174
rect 170288 114854 170608 114938
rect 170288 114618 170330 114854
rect 170566 114618 170608 114854
rect 170288 114586 170608 114618
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 168114 61774 168734 97218
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 168114 25774 168734 61218
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 101494 172454 136938
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 171834 65494 172454 100938
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 281537 186134 294618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 281537 189854 298338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 281537 193574 302058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 196674 594334 197294 629778
rect 196674 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 197294 594334
rect 196674 594014 197294 594098
rect 196674 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 197294 594014
rect 196674 558334 197294 593778
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 196674 486334 197294 521778
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 196674 450334 197294 485778
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 196674 414334 197294 449778
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 196674 378334 197294 413778
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 196674 281537 197294 305778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 598054 201014 633498
rect 200394 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 201014 598054
rect 200394 597734 201014 597818
rect 200394 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 201014 597734
rect 200394 562054 201014 597498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 601774 204734 637218
rect 204114 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 204734 601774
rect 204114 601454 204734 601538
rect 204114 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 204734 601454
rect 204114 565774 204734 601218
rect 204114 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 204734 565774
rect 204114 565454 204734 565538
rect 203379 565452 203445 565453
rect 203379 565388 203380 565452
rect 203444 565388 203445 565452
rect 203379 565387 203445 565388
rect 200394 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 201014 562054
rect 200394 561734 201014 561818
rect 200394 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 201014 561734
rect 200394 526054 201014 561498
rect 200394 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 201014 526054
rect 200394 525734 201014 525818
rect 200394 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 201014 525734
rect 200394 490054 201014 525498
rect 200394 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 201014 490054
rect 200394 489734 201014 489818
rect 200394 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 201014 489734
rect 200394 454054 201014 489498
rect 200394 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 201014 454054
rect 200394 453734 201014 453818
rect 200394 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 201014 453734
rect 200394 418054 201014 453498
rect 200394 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 201014 418054
rect 200394 417734 201014 417818
rect 200394 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 201014 417734
rect 200394 382054 201014 417498
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 281537 201014 309498
rect 203382 293317 203442 565387
rect 204114 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 204734 565454
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 214419 700772 214485 700773
rect 214419 700708 214420 700772
rect 214484 700708 214485 700772
rect 214419 700707 214485 700708
rect 211659 700636 211725 700637
rect 211659 700572 211660 700636
rect 211724 700572 211725 700636
rect 211659 700571 211725 700572
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 605494 208454 640938
rect 207834 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 208454 605494
rect 207834 605174 208454 605258
rect 207834 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 208454 605174
rect 207834 569494 208454 604938
rect 210739 596324 210805 596325
rect 210739 596260 210740 596324
rect 210804 596260 210805 596324
rect 210739 596259 210805 596260
rect 207834 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 208454 569494
rect 207834 569174 208454 569258
rect 207834 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 208454 569174
rect 206139 565316 206205 565317
rect 206139 565252 206140 565316
rect 206204 565252 206205 565316
rect 206139 565251 206205 565252
rect 204114 529774 204734 565218
rect 204114 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 204734 529774
rect 204114 529454 204734 529538
rect 204114 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 204734 529454
rect 204114 493774 204734 529218
rect 204114 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 204734 493774
rect 204114 493454 204734 493538
rect 204114 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 204734 493454
rect 204114 457774 204734 493218
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 204114 421774 204734 457218
rect 204114 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 204734 421774
rect 204114 421454 204734 421538
rect 204114 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 204734 421454
rect 204114 385774 204734 421218
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 203379 293316 203445 293317
rect 203379 293252 203380 293316
rect 203444 293252 203445 293316
rect 203379 293251 203445 293252
rect 204114 281537 204734 313218
rect 206142 293453 206202 565251
rect 206323 565180 206389 565181
rect 206323 565116 206324 565180
rect 206388 565116 206389 565180
rect 206323 565115 206389 565116
rect 206326 293589 206386 565115
rect 207834 533494 208454 568938
rect 208715 565044 208781 565045
rect 208715 564980 208716 565044
rect 208780 564980 208781 565044
rect 208715 564979 208781 564980
rect 207834 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 208454 533494
rect 207834 533174 208454 533258
rect 207834 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 208454 533174
rect 207834 497494 208454 532938
rect 207834 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 208454 497494
rect 207834 497174 208454 497258
rect 207834 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 208454 497174
rect 207834 461494 208454 496938
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 207834 425494 208454 460938
rect 207834 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 208454 425494
rect 207834 425174 208454 425258
rect 207834 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 208454 425174
rect 207834 389494 208454 424938
rect 207834 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 208454 389494
rect 207834 389174 208454 389258
rect 207834 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 208454 389174
rect 207834 353494 208454 388938
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 206323 293588 206389 293589
rect 206323 293524 206324 293588
rect 206388 293524 206389 293588
rect 206323 293523 206389 293524
rect 206139 293452 206205 293453
rect 206139 293388 206140 293452
rect 206204 293388 206205 293452
rect 206139 293387 206205 293388
rect 207834 281537 208454 316938
rect 208718 282845 208778 564979
rect 210742 358461 210802 596259
rect 210923 566540 210989 566541
rect 210923 566476 210924 566540
rect 210988 566476 210989 566540
rect 210923 566475 210989 566476
rect 210739 358460 210805 358461
rect 210739 358396 210740 358460
rect 210804 358396 210805 358460
rect 210739 358395 210805 358396
rect 210926 282845 210986 566475
rect 211662 342957 211722 700571
rect 213131 700364 213197 700365
rect 213131 700300 213132 700364
rect 213196 700300 213197 700364
rect 213131 700299 213197 700300
rect 212395 571980 212461 571981
rect 212395 571916 212396 571980
rect 212460 571916 212461 571980
rect 212395 571915 212461 571916
rect 212211 460188 212277 460189
rect 212211 460124 212212 460188
rect 212276 460124 212277 460188
rect 212211 460123 212277 460124
rect 211659 342956 211725 342957
rect 211659 342892 211660 342956
rect 211724 342892 211725 342956
rect 211659 342891 211725 342892
rect 212214 282845 212274 460123
rect 208715 282844 208781 282845
rect 208715 282780 208716 282844
rect 208780 282780 208781 282844
rect 208715 282779 208781 282780
rect 210923 282844 210989 282845
rect 210923 282780 210924 282844
rect 210988 282780 210989 282844
rect 210923 282779 210989 282780
rect 212211 282844 212277 282845
rect 212211 282780 212212 282844
rect 212276 282780 212277 282844
rect 212211 282779 212277 282780
rect 212398 282709 212458 571915
rect 212579 566404 212645 566405
rect 212579 566340 212580 566404
rect 212644 566340 212645 566404
rect 212579 566339 212645 566340
rect 212582 282709 212642 566339
rect 213134 337381 213194 700299
rect 213131 337380 213197 337381
rect 213131 337316 213132 337380
rect 213196 337316 213197 337380
rect 213131 337315 213197 337316
rect 214422 327725 214482 700707
rect 215891 700500 215957 700501
rect 215891 700436 215892 700500
rect 215956 700436 215957 700500
rect 215891 700435 215957 700436
rect 215155 594148 215221 594149
rect 215155 594084 215156 594148
rect 215220 594084 215221 594148
rect 215155 594083 215221 594084
rect 214787 445228 214853 445229
rect 214787 445164 214788 445228
rect 214852 445164 214853 445228
rect 214787 445163 214853 445164
rect 214603 445092 214669 445093
rect 214603 445028 214604 445092
rect 214668 445028 214669 445092
rect 214603 445027 214669 445028
rect 214419 327724 214485 327725
rect 214419 327660 214420 327724
rect 214484 327660 214485 327724
rect 214419 327659 214485 327660
rect 214606 287877 214666 445027
rect 214603 287876 214669 287877
rect 214603 287812 214604 287876
rect 214668 287812 214669 287876
rect 214603 287811 214669 287812
rect 214790 287741 214850 445163
rect 215158 355469 215218 594083
rect 215155 355468 215221 355469
rect 215155 355404 215156 355468
rect 215220 355404 215221 355468
rect 215155 355403 215221 355404
rect 215894 355333 215954 700435
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 685244 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 685244 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 685244 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 685244 229574 698058
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 685244 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 685244 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 685244 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 685244 265574 698058
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 685244 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 685244 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 685244 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 685244 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 685244 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 685244 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 685244 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 685244 337574 698058
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 350947 685948 351013 685949
rect 350947 685884 350948 685948
rect 351012 685884 351013 685948
rect 350947 685883 351013 685884
rect 350950 683770 351010 685883
rect 350840 683710 351010 683770
rect 350840 683202 350900 683710
rect 220272 655174 220620 655206
rect 220272 654938 220328 655174
rect 220564 654938 220620 655174
rect 220272 654854 220620 654938
rect 220272 654618 220328 654854
rect 220564 654618 220620 654854
rect 220272 654586 220620 654618
rect 356000 655174 356348 655206
rect 356000 654938 356056 655174
rect 356292 654938 356348 655174
rect 356000 654854 356348 654938
rect 356000 654618 356056 654854
rect 356292 654618 356348 654854
rect 356000 654586 356348 654618
rect 220952 651454 221300 651486
rect 220952 651218 221008 651454
rect 221244 651218 221300 651454
rect 220952 651134 221300 651218
rect 220952 650898 221008 651134
rect 221244 650898 221300 651134
rect 220952 650866 221300 650898
rect 355320 651454 355668 651486
rect 355320 651218 355376 651454
rect 355612 651218 355668 651454
rect 355320 651134 355668 651218
rect 355320 650898 355376 651134
rect 355612 650898 355668 651134
rect 355320 650866 355668 650898
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 220272 619174 220620 619206
rect 220272 618938 220328 619174
rect 220564 618938 220620 619174
rect 220272 618854 220620 618938
rect 220272 618618 220328 618854
rect 220564 618618 220620 618854
rect 220272 618586 220620 618618
rect 356000 619174 356348 619206
rect 356000 618938 356056 619174
rect 356292 618938 356348 619174
rect 356000 618854 356348 618938
rect 356000 618618 356056 618854
rect 356292 618618 356348 618854
rect 356000 618586 356348 618618
rect 220952 615454 221300 615486
rect 220952 615218 221008 615454
rect 221244 615218 221300 615454
rect 220952 615134 221300 615218
rect 220952 614898 221008 615134
rect 221244 614898 221300 615134
rect 220952 614866 221300 614898
rect 355320 615454 355668 615486
rect 355320 615218 355376 615454
rect 355612 615218 355668 615454
rect 355320 615134 355668 615218
rect 355320 614898 355376 615134
rect 355612 614898 355668 615134
rect 355320 614866 355668 614898
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 219203 608020 219269 608021
rect 219203 607956 219204 608020
rect 219268 607956 219269 608020
rect 219203 607955 219269 607956
rect 219019 597276 219085 597277
rect 219019 597212 219020 597276
rect 219084 597212 219085 597276
rect 219019 597211 219085 597212
rect 216259 596596 216325 596597
rect 216259 596532 216260 596596
rect 216324 596532 216325 596596
rect 216259 596531 216325 596532
rect 216075 461548 216141 461549
rect 216075 461484 216076 461548
rect 216140 461484 216141 461548
rect 216075 461483 216141 461484
rect 215891 355332 215957 355333
rect 215891 355268 215892 355332
rect 215956 355268 215957 355332
rect 215891 355267 215957 355268
rect 214787 287740 214853 287741
rect 214787 287676 214788 287740
rect 214852 287676 214853 287740
rect 214787 287675 214853 287676
rect 216078 282845 216138 461483
rect 216262 358733 216322 596531
rect 217731 594012 217797 594013
rect 217731 593948 217732 594012
rect 217796 593948 217797 594012
rect 217731 593947 217797 593948
rect 216443 570620 216509 570621
rect 216443 570556 216444 570620
rect 216508 570556 216509 570620
rect 216443 570555 216509 570556
rect 216259 358732 216325 358733
rect 216259 358668 216260 358732
rect 216324 358668 216325 358732
rect 216259 358667 216325 358668
rect 216446 282845 216506 570555
rect 217179 478956 217245 478957
rect 217179 478892 217180 478956
rect 217244 478892 217245 478956
rect 217179 478891 217245 478892
rect 216811 444956 216877 444957
rect 216811 444892 216812 444956
rect 216876 444892 216877 444956
rect 216811 444891 216877 444892
rect 216627 443596 216693 443597
rect 216627 443532 216628 443596
rect 216692 443532 216693 443596
rect 216627 443531 216693 443532
rect 216630 282845 216690 443531
rect 216814 369885 216874 444891
rect 217182 393821 217242 478891
rect 217734 474741 217794 593947
rect 218651 570756 218717 570757
rect 218651 570692 218652 570756
rect 218716 570692 218717 570756
rect 218651 570691 218717 570692
rect 217915 567220 217981 567221
rect 217915 567156 217916 567220
rect 217980 567156 217981 567220
rect 217915 567155 217981 567156
rect 217918 488341 217978 567155
rect 217915 488340 217981 488341
rect 217915 488276 217916 488340
rect 217980 488276 217981 488340
rect 217915 488275 217981 488276
rect 217918 487253 217978 488275
rect 217915 487252 217981 487253
rect 217915 487188 217916 487252
rect 217980 487188 217981 487252
rect 217915 487187 217981 487188
rect 217731 474740 217797 474741
rect 217731 474676 217732 474740
rect 217796 474676 217797 474740
rect 217731 474675 217797 474676
rect 217731 393956 217797 393957
rect 217731 393892 217732 393956
rect 217796 393892 217797 393956
rect 217731 393891 217797 393892
rect 217179 393820 217245 393821
rect 217179 393756 217180 393820
rect 217244 393756 217245 393820
rect 217179 393755 217245 393756
rect 217363 370020 217429 370021
rect 217363 369956 217364 370020
rect 217428 369956 217429 370020
rect 217363 369955 217429 369956
rect 216811 369884 216877 369885
rect 216811 369820 216812 369884
rect 216876 369820 216877 369884
rect 216811 369819 216877 369820
rect 217366 342957 217426 369955
rect 217547 368388 217613 368389
rect 217547 368324 217548 368388
rect 217612 368324 217613 368388
rect 217547 368323 217613 368324
rect 217363 342956 217429 342957
rect 217363 342892 217364 342956
rect 217428 342892 217429 342956
rect 217363 342891 217429 342892
rect 216075 282844 216141 282845
rect 216075 282780 216076 282844
rect 216140 282780 216141 282844
rect 216075 282779 216141 282780
rect 216443 282844 216509 282845
rect 216443 282780 216444 282844
rect 216508 282780 216509 282844
rect 216443 282779 216509 282780
rect 216627 282844 216693 282845
rect 216627 282780 216628 282844
rect 216692 282780 216693 282844
rect 216627 282779 216693 282780
rect 212395 282708 212461 282709
rect 212395 282644 212396 282708
rect 212460 282644 212461 282708
rect 212395 282643 212461 282644
rect 212579 282708 212645 282709
rect 212579 282644 212580 282708
rect 212644 282644 212645 282708
rect 212579 282643 212645 282644
rect 217550 282573 217610 368323
rect 217734 359685 217794 393891
rect 217918 368389 217978 487187
rect 217915 368388 217981 368389
rect 217915 368324 217916 368388
rect 217980 368324 217981 368388
rect 217915 368323 217981 368324
rect 217731 359684 217797 359685
rect 217731 359620 217732 359684
rect 217796 359620 217797 359684
rect 217731 359619 217797 359620
rect 217794 327454 218414 358064
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217547 282572 217613 282573
rect 217547 282508 217548 282572
rect 217612 282508 217613 282572
rect 217547 282507 217613 282508
rect 217794 281537 218414 290898
rect 218654 282845 218714 570691
rect 218835 474740 218901 474741
rect 218835 474676 218836 474740
rect 218900 474676 218901 474740
rect 218835 474675 218901 474676
rect 218838 359413 218898 474675
rect 218835 359412 218901 359413
rect 218835 359348 218836 359412
rect 218900 359348 218901 359412
rect 218835 359347 218901 359348
rect 219022 358189 219082 597211
rect 219206 359957 219266 607955
rect 357939 607476 358005 607477
rect 357939 607412 357940 607476
rect 358004 607412 358005 607476
rect 357939 607411 358005 607412
rect 236056 599450 236116 600100
rect 237144 599450 237204 600100
rect 238232 599450 238292 600100
rect 239592 599586 239652 600100
rect 238894 599526 239652 599586
rect 240544 599586 240604 600100
rect 241768 599586 241828 600100
rect 243128 599586 243188 600100
rect 240544 599526 240610 599586
rect 238894 599450 238954 599526
rect 235950 599390 236116 599450
rect 237054 599390 237204 599450
rect 238158 599390 238292 599450
rect 238526 599390 238954 599450
rect 235950 597549 236010 599390
rect 237054 597549 237114 599390
rect 238158 597549 238218 599390
rect 235947 597548 236013 597549
rect 235947 597484 235948 597548
rect 236012 597484 236013 597548
rect 235947 597483 236013 597484
rect 237051 597548 237117 597549
rect 237051 597484 237052 597548
rect 237116 597484 237117 597548
rect 237051 597483 237117 597484
rect 238155 597548 238221 597549
rect 238155 597484 238156 597548
rect 238220 597484 238221 597548
rect 238155 597483 238221 597484
rect 238526 596869 238586 599390
rect 240550 596869 240610 599526
rect 241654 599526 241828 599586
rect 243126 599526 243188 599586
rect 244216 599586 244276 600100
rect 245440 599586 245500 600100
rect 246528 599586 246588 600100
rect 247616 599586 247676 600100
rect 248296 599586 248356 600100
rect 248704 599586 248764 600100
rect 244216 599526 244290 599586
rect 245440 599526 245578 599586
rect 241654 596869 241714 599526
rect 243126 597549 243186 599526
rect 244230 597549 244290 599526
rect 245518 597549 245578 599526
rect 246438 599526 246588 599586
rect 247542 599526 247676 599586
rect 248278 599526 248356 599586
rect 248646 599526 248764 599586
rect 250064 599586 250124 600100
rect 250744 599586 250804 600100
rect 250064 599526 250178 599586
rect 246438 597549 246498 599526
rect 243123 597548 243189 597549
rect 243123 597484 243124 597548
rect 243188 597484 243189 597548
rect 243123 597483 243189 597484
rect 244227 597548 244293 597549
rect 244227 597484 244228 597548
rect 244292 597484 244293 597548
rect 244227 597483 244293 597484
rect 245515 597548 245581 597549
rect 245515 597484 245516 597548
rect 245580 597484 245581 597548
rect 245515 597483 245581 597484
rect 246435 597548 246501 597549
rect 246435 597484 246436 597548
rect 246500 597484 246501 597548
rect 246435 597483 246501 597484
rect 247542 596869 247602 599526
rect 248278 597549 248338 599526
rect 248646 597549 248706 599526
rect 248275 597548 248341 597549
rect 248275 597484 248276 597548
rect 248340 597484 248341 597548
rect 248275 597483 248341 597484
rect 248643 597548 248709 597549
rect 248643 597484 248644 597548
rect 248708 597484 248709 597548
rect 248643 597483 248709 597484
rect 250118 596869 250178 599526
rect 250670 599526 250804 599586
rect 251288 599586 251348 600100
rect 252376 599586 252436 600100
rect 253464 599586 253524 600100
rect 251288 599526 251466 599586
rect 250670 597549 250730 599526
rect 250667 597548 250733 597549
rect 250667 597484 250668 597548
rect 250732 597484 250733 597548
rect 250667 597483 250733 597484
rect 251406 596869 251466 599526
rect 252326 599526 252436 599586
rect 253430 599526 253524 599586
rect 253600 599586 253660 600100
rect 254552 599586 254612 600100
rect 255912 599586 255972 600100
rect 253600 599526 253674 599586
rect 252326 597549 252386 599526
rect 253430 597549 253490 599526
rect 252323 597548 252389 597549
rect 252323 597484 252324 597548
rect 252388 597484 252389 597548
rect 252323 597483 252389 597484
rect 253427 597548 253493 597549
rect 253427 597484 253428 597548
rect 253492 597484 253493 597548
rect 253427 597483 253493 597484
rect 219939 596868 220005 596869
rect 219939 596804 219940 596868
rect 220004 596804 220005 596868
rect 219939 596803 220005 596804
rect 238523 596868 238589 596869
rect 238523 596804 238524 596868
rect 238588 596804 238589 596868
rect 238523 596803 238589 596804
rect 240547 596868 240613 596869
rect 240547 596804 240548 596868
rect 240612 596804 240613 596868
rect 240547 596803 240613 596804
rect 241651 596868 241717 596869
rect 241651 596804 241652 596868
rect 241716 596804 241717 596868
rect 241651 596803 241717 596804
rect 247539 596868 247605 596869
rect 247539 596804 247540 596868
rect 247604 596804 247605 596868
rect 247539 596803 247605 596804
rect 250115 596868 250181 596869
rect 250115 596804 250116 596868
rect 250180 596804 250181 596868
rect 250115 596803 250181 596804
rect 251403 596868 251469 596869
rect 251403 596804 251404 596868
rect 251468 596804 251469 596868
rect 251403 596803 251469 596804
rect 219755 563684 219821 563685
rect 219755 563620 219756 563684
rect 219820 563620 219821 563684
rect 219755 563619 219821 563620
rect 219203 359956 219269 359957
rect 219203 359892 219204 359956
rect 219268 359892 219269 359956
rect 219203 359891 219269 359892
rect 219019 358188 219085 358189
rect 219019 358124 219020 358188
rect 219084 358124 219085 358188
rect 219019 358123 219085 358124
rect 219758 282845 219818 563619
rect 219942 289101 220002 596803
rect 253614 596325 253674 599526
rect 254534 599526 254612 599586
rect 255822 599526 255972 599586
rect 254534 597549 254594 599526
rect 255822 597549 255882 599526
rect 256048 599450 256108 600100
rect 257000 599586 257060 600100
rect 258088 599589 258148 600100
rect 256006 599390 256108 599450
rect 256926 599526 257060 599586
rect 258085 599588 258151 599589
rect 254531 597548 254597 597549
rect 254531 597484 254532 597548
rect 254596 597484 254597 597548
rect 254531 597483 254597 597484
rect 255819 597548 255885 597549
rect 255819 597484 255820 597548
rect 255884 597484 255885 597548
rect 255819 597483 255885 597484
rect 256006 596597 256066 599390
rect 256926 597549 256986 599526
rect 258085 599524 258086 599588
rect 258150 599524 258151 599588
rect 258085 599523 258151 599524
rect 258496 599450 258556 600100
rect 258214 599390 258556 599450
rect 259448 599450 259508 600100
rect 260672 599450 260732 600100
rect 261080 599450 261140 600100
rect 261760 599450 261820 600100
rect 262848 599450 262908 600100
rect 259448 599390 259562 599450
rect 258214 598950 258274 599390
rect 257846 598890 258274 598950
rect 256923 597548 256989 597549
rect 256923 597484 256924 597548
rect 256988 597484 256989 597548
rect 256923 597483 256989 597484
rect 257846 596733 257906 598890
rect 259502 596733 259562 599390
rect 260606 599390 260732 599450
rect 260974 599390 261140 599450
rect 261710 599390 261820 599450
rect 262814 599390 262908 599450
rect 263528 599450 263588 600100
rect 263936 599450 263996 600100
rect 265296 599450 265356 600100
rect 265976 599450 266036 600100
rect 266384 599450 266444 600100
rect 267608 599450 267668 600100
rect 268288 599586 268348 600100
rect 268696 599586 268756 600100
rect 269784 599586 269844 600100
rect 271008 599586 271068 600100
rect 268288 599526 268394 599586
rect 268696 599526 268762 599586
rect 269784 599526 269866 599586
rect 263528 599390 263610 599450
rect 257843 596732 257909 596733
rect 257843 596668 257844 596732
rect 257908 596668 257909 596732
rect 257843 596667 257909 596668
rect 259499 596732 259565 596733
rect 259499 596668 259500 596732
rect 259564 596668 259565 596732
rect 259499 596667 259565 596668
rect 260606 596597 260666 599390
rect 260974 597413 261034 599390
rect 261710 597549 261770 599390
rect 261707 597548 261773 597549
rect 261707 597484 261708 597548
rect 261772 597484 261773 597548
rect 261707 597483 261773 597484
rect 262814 597413 262874 599390
rect 263550 597549 263610 599390
rect 263918 599390 263996 599450
rect 265206 599390 265356 599450
rect 265942 599390 266036 599450
rect 266310 599390 266444 599450
rect 267598 599390 267668 599450
rect 263547 597548 263613 597549
rect 263547 597484 263548 597548
rect 263612 597484 263613 597548
rect 263547 597483 263613 597484
rect 263918 597413 263978 599390
rect 260971 597412 261037 597413
rect 260971 597348 260972 597412
rect 261036 597348 261037 597412
rect 260971 597347 261037 597348
rect 262811 597412 262877 597413
rect 262811 597348 262812 597412
rect 262876 597348 262877 597412
rect 262811 597347 262877 597348
rect 263915 597412 263981 597413
rect 263915 597348 263916 597412
rect 263980 597348 263981 597412
rect 263915 597347 263981 597348
rect 265206 596869 265266 599390
rect 265942 597549 266002 599390
rect 265939 597548 266005 597549
rect 265939 597484 265940 597548
rect 266004 597484 266005 597548
rect 265939 597483 266005 597484
rect 265203 596868 265269 596869
rect 265203 596804 265204 596868
rect 265268 596804 265269 596868
rect 265203 596803 265269 596804
rect 256003 596596 256069 596597
rect 256003 596532 256004 596596
rect 256068 596532 256069 596596
rect 256003 596531 256069 596532
rect 260603 596596 260669 596597
rect 260603 596532 260604 596596
rect 260668 596532 260669 596596
rect 260603 596531 260669 596532
rect 266310 596461 266370 599390
rect 267598 597413 267658 599390
rect 268334 597549 268394 599526
rect 268331 597548 268397 597549
rect 268331 597484 268332 597548
rect 268396 597484 268397 597548
rect 268331 597483 268397 597484
rect 267595 597412 267661 597413
rect 267595 597348 267596 597412
rect 267660 597348 267661 597412
rect 267595 597347 267661 597348
rect 268702 596733 268762 599526
rect 269806 596733 269866 599526
rect 270910 599526 271068 599586
rect 270910 597549 270970 599526
rect 271144 599450 271204 600100
rect 272232 599586 272292 600100
rect 273320 599586 273380 600100
rect 273592 599586 273652 600100
rect 274408 599586 274468 600100
rect 275768 599586 275828 600100
rect 271094 599390 271204 599450
rect 272198 599526 272292 599586
rect 273302 599526 273380 599586
rect 273486 599526 273652 599586
rect 274406 599526 274468 599586
rect 275694 599526 275828 599586
rect 276040 599586 276100 600100
rect 276992 599586 277052 600100
rect 276040 599526 276122 599586
rect 270907 597548 270973 597549
rect 270907 597484 270908 597548
rect 270972 597484 270973 597548
rect 270907 597483 270973 597484
rect 271094 597141 271154 599390
rect 271091 597140 271157 597141
rect 271091 597076 271092 597140
rect 271156 597076 271157 597140
rect 271091 597075 271157 597076
rect 268699 596732 268765 596733
rect 268699 596668 268700 596732
rect 268764 596668 268765 596732
rect 268699 596667 268765 596668
rect 269803 596732 269869 596733
rect 269803 596668 269804 596732
rect 269868 596668 269869 596732
rect 269803 596667 269869 596668
rect 272198 596461 272258 599526
rect 273302 597141 273362 599526
rect 273486 597277 273546 599526
rect 273483 597276 273549 597277
rect 273483 597212 273484 597276
rect 273548 597212 273549 597276
rect 273483 597211 273549 597212
rect 273299 597140 273365 597141
rect 273299 597076 273300 597140
rect 273364 597076 273365 597140
rect 273299 597075 273365 597076
rect 266307 596460 266373 596461
rect 266307 596396 266308 596460
rect 266372 596396 266373 596460
rect 266307 596395 266373 596396
rect 272195 596460 272261 596461
rect 272195 596396 272196 596460
rect 272260 596396 272261 596460
rect 272195 596395 272261 596396
rect 274406 596325 274466 599526
rect 275694 597277 275754 599526
rect 276062 597413 276122 599526
rect 276982 599526 277052 599586
rect 278080 599586 278140 600100
rect 278488 599589 278548 600100
rect 278485 599588 278551 599589
rect 278080 599526 278146 599586
rect 276982 597549 277042 599526
rect 276979 597548 277045 597549
rect 276979 597484 276980 597548
rect 277044 597484 277045 597548
rect 276979 597483 277045 597484
rect 276059 597412 276125 597413
rect 276059 597348 276060 597412
rect 276124 597348 276125 597412
rect 276059 597347 276125 597348
rect 275691 597276 275757 597277
rect 275691 597212 275692 597276
rect 275756 597212 275757 597276
rect 275691 597211 275757 597212
rect 278086 596869 278146 599526
rect 278485 599524 278486 599588
rect 278550 599524 278551 599588
rect 279168 599586 279228 600100
rect 280936 599586 280996 600100
rect 283520 599586 283580 600100
rect 279168 599526 279250 599586
rect 278485 599523 278551 599524
rect 278083 596868 278149 596869
rect 278083 596804 278084 596868
rect 278148 596804 278149 596868
rect 278083 596803 278149 596804
rect 279190 596597 279250 599526
rect 280846 599526 280996 599586
rect 283422 599526 283580 599586
rect 285968 599586 286028 600100
rect 285968 599526 286058 599586
rect 280846 597549 280906 599526
rect 283422 597549 283482 599526
rect 285998 597549 286058 599526
rect 288280 599450 288340 600100
rect 291000 599450 291060 600100
rect 293448 599450 293508 600100
rect 288206 599390 288340 599450
rect 290966 599390 291060 599450
rect 293358 599390 293508 599450
rect 295896 599450 295956 600100
rect 298480 599450 298540 600100
rect 300928 599450 300988 600100
rect 303512 599450 303572 600100
rect 295896 599390 295994 599450
rect 298480 599390 298570 599450
rect 280843 597548 280909 597549
rect 280843 597484 280844 597548
rect 280908 597484 280909 597548
rect 280843 597483 280909 597484
rect 283419 597548 283485 597549
rect 283419 597484 283420 597548
rect 283484 597484 283485 597548
rect 283419 597483 283485 597484
rect 285995 597548 286061 597549
rect 285995 597484 285996 597548
rect 286060 597484 286061 597548
rect 285995 597483 286061 597484
rect 288206 597141 288266 599390
rect 290966 597549 291026 599390
rect 293358 597549 293418 599390
rect 290963 597548 291029 597549
rect 290963 597484 290964 597548
rect 291028 597484 291029 597548
rect 290963 597483 291029 597484
rect 293355 597548 293421 597549
rect 293355 597484 293356 597548
rect 293420 597484 293421 597548
rect 293355 597483 293421 597484
rect 288203 597140 288269 597141
rect 288203 597076 288204 597140
rect 288268 597076 288269 597140
rect 288203 597075 288269 597076
rect 279187 596596 279253 596597
rect 279187 596532 279188 596596
rect 279252 596532 279253 596596
rect 279187 596531 279253 596532
rect 295934 596325 295994 599390
rect 298510 597277 298570 599390
rect 300902 599390 300988 599450
rect 303478 599390 303572 599450
rect 305960 599450 306020 600100
rect 308544 599450 308604 600100
rect 310992 599450 311052 600100
rect 313440 599450 313500 600100
rect 315888 599450 315948 600100
rect 305960 599390 306114 599450
rect 308544 599390 308690 599450
rect 310992 599390 311082 599450
rect 300902 597413 300962 599390
rect 300899 597412 300965 597413
rect 300899 597348 300900 597412
rect 300964 597348 300965 597412
rect 300899 597347 300965 597348
rect 298507 597276 298573 597277
rect 298507 597212 298508 597276
rect 298572 597212 298573 597276
rect 298507 597211 298573 597212
rect 303478 596325 303538 599390
rect 306054 596461 306114 599390
rect 308630 596461 308690 599390
rect 311022 596869 311082 599390
rect 313414 599390 313500 599450
rect 315806 599390 315948 599450
rect 318472 599450 318532 600100
rect 320920 599450 320980 600100
rect 323368 599450 323428 600100
rect 325952 599450 326012 600100
rect 318472 599390 318626 599450
rect 320920 599390 321018 599450
rect 311019 596868 311085 596869
rect 311019 596804 311020 596868
rect 311084 596804 311085 596868
rect 311019 596803 311085 596804
rect 313414 596733 313474 599390
rect 313411 596732 313477 596733
rect 313411 596668 313412 596732
rect 313476 596668 313477 596732
rect 313411 596667 313477 596668
rect 315806 596597 315866 599390
rect 318566 596733 318626 599390
rect 320958 596869 321018 599390
rect 323350 599390 323428 599450
rect 325926 599390 326012 599450
rect 323350 596869 323410 599390
rect 325926 597005 325986 599390
rect 357571 597412 357637 597413
rect 357571 597348 357572 597412
rect 357636 597348 357637 597412
rect 357571 597347 357637 597348
rect 357019 597140 357085 597141
rect 357019 597076 357020 597140
rect 357084 597076 357085 597140
rect 357019 597075 357085 597076
rect 325923 597004 325989 597005
rect 325923 596940 325924 597004
rect 325988 596940 325989 597004
rect 325923 596939 325989 596940
rect 356651 597004 356717 597005
rect 356651 596940 356652 597004
rect 356716 596940 356717 597004
rect 356651 596939 356717 596940
rect 320955 596868 321021 596869
rect 320955 596804 320956 596868
rect 321020 596804 321021 596868
rect 320955 596803 321021 596804
rect 323347 596868 323413 596869
rect 323347 596804 323348 596868
rect 323412 596804 323413 596868
rect 323347 596803 323413 596804
rect 318563 596732 318629 596733
rect 318563 596668 318564 596732
rect 318628 596668 318629 596732
rect 318563 596667 318629 596668
rect 315803 596596 315869 596597
rect 315803 596532 315804 596596
rect 315868 596532 315869 596596
rect 315803 596531 315869 596532
rect 306051 596460 306117 596461
rect 306051 596396 306052 596460
rect 306116 596396 306117 596460
rect 306051 596395 306117 596396
rect 308627 596460 308693 596461
rect 308627 596396 308628 596460
rect 308692 596396 308693 596460
rect 308627 596395 308693 596396
rect 253611 596324 253677 596325
rect 253611 596260 253612 596324
rect 253676 596260 253677 596324
rect 253611 596259 253677 596260
rect 274403 596324 274469 596325
rect 274403 596260 274404 596324
rect 274468 596260 274469 596324
rect 274403 596259 274469 596260
rect 295931 596324 295997 596325
rect 295931 596260 295932 596324
rect 295996 596260 295997 596324
rect 295931 596259 295997 596260
rect 303475 596324 303541 596325
rect 303475 596260 303476 596324
rect 303540 596260 303541 596324
rect 303475 596259 303541 596260
rect 350947 565860 351013 565861
rect 350947 565796 350948 565860
rect 351012 565796 351013 565860
rect 350947 565795 351013 565796
rect 350950 564090 351010 565795
rect 350840 564030 351010 564090
rect 350840 563202 350900 564030
rect 220272 547174 220620 547206
rect 220272 546938 220328 547174
rect 220564 546938 220620 547174
rect 220272 546854 220620 546938
rect 220272 546618 220328 546854
rect 220564 546618 220620 546854
rect 220272 546586 220620 546618
rect 356000 547174 356348 547206
rect 356000 546938 356056 547174
rect 356292 546938 356348 547174
rect 356000 546854 356348 546938
rect 356000 546618 356056 546854
rect 356292 546618 356348 546854
rect 356000 546586 356348 546618
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 220272 511174 220620 511206
rect 220272 510938 220328 511174
rect 220564 510938 220620 511174
rect 220272 510854 220620 510938
rect 220272 510618 220328 510854
rect 220564 510618 220620 510854
rect 220272 510586 220620 510618
rect 356000 511174 356348 511206
rect 356000 510938 356056 511174
rect 356292 510938 356348 511174
rect 356000 510854 356348 510938
rect 356000 510618 356056 510854
rect 356292 510618 356348 510854
rect 356000 510586 356348 510618
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 236056 479637 236116 480080
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 237054 479710 237204 479770
rect 238158 479710 238292 479770
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 236053 479636 236119 479637
rect 236053 479572 236054 479636
rect 236118 479572 236119 479636
rect 236053 479571 236119 479572
rect 237054 477325 237114 479710
rect 237051 477324 237117 477325
rect 237051 477260 237052 477324
rect 237116 477260 237117 477324
rect 237051 477259 237117 477260
rect 238158 476917 238218 479710
rect 239630 477461 239690 479710
rect 239627 477460 239693 477461
rect 239627 477396 239628 477460
rect 239692 477396 239693 477460
rect 239627 477395 239693 477396
rect 240550 477053 240610 479710
rect 241654 479710 241828 479770
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 245440 479710 245578 479770
rect 241654 477189 241714 479710
rect 243126 477461 243186 479710
rect 244230 477461 244290 479710
rect 245518 477461 245578 479710
rect 246438 479710 246588 479770
rect 247542 479710 247676 479770
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 250064 479710 250178 479770
rect 246438 477461 246498 479710
rect 247542 477461 247602 479710
rect 243123 477460 243189 477461
rect 243123 477396 243124 477460
rect 243188 477396 243189 477460
rect 243123 477395 243189 477396
rect 244227 477460 244293 477461
rect 244227 477396 244228 477460
rect 244292 477396 244293 477460
rect 244227 477395 244293 477396
rect 245515 477460 245581 477461
rect 245515 477396 245516 477460
rect 245580 477396 245581 477460
rect 245515 477395 245581 477396
rect 246435 477460 246501 477461
rect 246435 477396 246436 477460
rect 246500 477396 246501 477460
rect 246435 477395 246501 477396
rect 247539 477460 247605 477461
rect 247539 477396 247540 477460
rect 247604 477396 247605 477460
rect 247539 477395 247605 477396
rect 241651 477188 241717 477189
rect 241651 477124 241652 477188
rect 241716 477124 241717 477188
rect 241651 477123 241717 477124
rect 240547 477052 240613 477053
rect 240547 476988 240548 477052
rect 240612 476988 240613 477052
rect 240547 476987 240613 476988
rect 238155 476916 238221 476917
rect 238155 476852 238156 476916
rect 238220 476852 238221 476916
rect 238155 476851 238221 476852
rect 248278 476237 248338 479710
rect 248646 477461 248706 479710
rect 250118 477461 250178 479710
rect 250670 479710 250804 479770
rect 251222 479710 251348 479770
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 248643 477460 248709 477461
rect 248643 477396 248644 477460
rect 248708 477396 248709 477460
rect 248643 477395 248709 477396
rect 250115 477460 250181 477461
rect 250115 477396 250116 477460
rect 250180 477396 250181 477460
rect 250115 477395 250181 477396
rect 250670 476237 250730 479710
rect 251222 477461 251282 479710
rect 252326 477461 252386 479710
rect 253430 477461 253490 479710
rect 251219 477460 251285 477461
rect 251219 477396 251220 477460
rect 251284 477396 251285 477460
rect 251219 477395 251285 477396
rect 252323 477460 252389 477461
rect 252323 477396 252324 477460
rect 252388 477396 252389 477460
rect 252323 477395 252389 477396
rect 253427 477460 253493 477461
rect 253427 477396 253428 477460
rect 253492 477396 253493 477460
rect 253427 477395 253493 477396
rect 253614 476237 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 258496 479770 258556 480080
rect 256048 479710 256250 479770
rect 254534 477461 254594 479710
rect 255822 477461 255882 479710
rect 254531 477460 254597 477461
rect 254531 477396 254532 477460
rect 254596 477396 254597 477460
rect 254531 477395 254597 477396
rect 255819 477460 255885 477461
rect 255819 477396 255820 477460
rect 255884 477396 255885 477460
rect 255819 477395 255885 477396
rect 256190 476917 256250 479710
rect 256926 479710 257060 479770
rect 257846 479710 258148 479770
rect 258398 479710 258556 479770
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 259448 479710 259562 479770
rect 260672 479710 260850 479770
rect 256926 477461 256986 479710
rect 257846 477730 257906 479710
rect 257846 477670 258274 477730
rect 256923 477460 256989 477461
rect 256923 477396 256924 477460
rect 256988 477396 256989 477460
rect 256923 477395 256989 477396
rect 258214 477325 258274 477670
rect 258211 477324 258277 477325
rect 258211 477260 258212 477324
rect 258276 477260 258277 477324
rect 258211 477259 258277 477260
rect 256187 476916 256253 476917
rect 256187 476852 256188 476916
rect 256252 476852 256253 476916
rect 256187 476851 256253 476852
rect 258398 476237 258458 479710
rect 259502 476645 259562 479710
rect 260790 477461 260850 479710
rect 260974 479710 261140 479770
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 263528 479710 263610 479770
rect 260787 477460 260853 477461
rect 260787 477396 260788 477460
rect 260852 477396 260853 477460
rect 260787 477395 260853 477396
rect 259499 476644 259565 476645
rect 259499 476580 259500 476644
rect 259564 476580 259565 476644
rect 259499 476579 259565 476580
rect 260790 476509 260850 477395
rect 260787 476508 260853 476509
rect 260787 476444 260788 476508
rect 260852 476444 260853 476508
rect 260787 476443 260853 476444
rect 260974 476237 261034 479710
rect 261710 477325 261770 479710
rect 261707 477324 261773 477325
rect 261707 477260 261708 477324
rect 261772 477260 261773 477324
rect 261707 477259 261773 477260
rect 262814 476917 262874 479710
rect 262811 476916 262877 476917
rect 262811 476852 262812 476916
rect 262876 476852 262877 476916
rect 262811 476851 262877 476852
rect 263550 476237 263610 479710
rect 263918 479710 263996 479770
rect 265206 479710 265356 479770
rect 265942 479710 266036 479770
rect 266310 479710 266444 479770
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 263918 477325 263978 479710
rect 263915 477324 263981 477325
rect 263915 477260 263916 477324
rect 263980 477260 263981 477324
rect 263915 477259 263981 477260
rect 265206 477053 265266 479710
rect 265203 477052 265269 477053
rect 265203 476988 265204 477052
rect 265268 476988 265269 477052
rect 265203 476987 265269 476988
rect 265942 476237 266002 479710
rect 266310 477461 266370 479710
rect 266307 477460 266373 477461
rect 266307 477396 266308 477460
rect 266372 477396 266373 477460
rect 266307 477395 266373 477396
rect 267598 476781 267658 479710
rect 267595 476780 267661 476781
rect 267595 476716 267596 476780
rect 267660 476716 267661 476780
rect 267595 476715 267661 476716
rect 268334 476237 268394 479710
rect 268702 476645 268762 479710
rect 269806 477461 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 275768 479770 275828 480080
rect 271144 479710 271338 479770
rect 269803 477460 269869 477461
rect 269803 477396 269804 477460
rect 269868 477396 269869 477460
rect 269803 477395 269869 477396
rect 270910 476917 270970 479710
rect 271278 477053 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273486 479710 273652 479770
rect 274406 479710 274468 479770
rect 275694 479710 275828 479770
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 276040 479710 276122 479770
rect 272198 477325 272258 479710
rect 272195 477324 272261 477325
rect 272195 477260 272196 477324
rect 272260 477260 272261 477324
rect 272195 477259 272261 477260
rect 271275 477052 271341 477053
rect 271275 476988 271276 477052
rect 271340 476988 271341 477052
rect 271275 476987 271341 476988
rect 273302 476917 273362 479710
rect 270907 476916 270973 476917
rect 270907 476852 270908 476916
rect 270972 476852 270973 476916
rect 270907 476851 270973 476852
rect 273299 476916 273365 476917
rect 273299 476852 273300 476916
rect 273364 476852 273365 476916
rect 273299 476851 273365 476852
rect 268699 476644 268765 476645
rect 268699 476580 268700 476644
rect 268764 476580 268765 476644
rect 268699 476579 268765 476580
rect 273486 476237 273546 479710
rect 274406 477189 274466 479710
rect 275694 477189 275754 479710
rect 274403 477188 274469 477189
rect 274403 477124 274404 477188
rect 274468 477124 274469 477188
rect 274403 477123 274469 477124
rect 275691 477188 275757 477189
rect 275691 477124 275692 477188
rect 275756 477124 275757 477188
rect 275691 477123 275757 477124
rect 276062 476237 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276982 477325 277042 479710
rect 278086 477325 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 279168 479710 279250 479770
rect 276979 477324 277045 477325
rect 276979 477260 276980 477324
rect 277044 477260 277045 477324
rect 276979 477259 277045 477260
rect 278083 477324 278149 477325
rect 278083 477260 278084 477324
rect 278148 477260 278149 477324
rect 278083 477259 278149 477260
rect 278454 477053 278514 479710
rect 279190 477461 279250 479710
rect 280846 479710 280996 479770
rect 283422 479710 283580 479770
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 293448 479770 293508 480080
rect 285968 479710 286058 479770
rect 279187 477460 279253 477461
rect 279187 477396 279188 477460
rect 279252 477396 279253 477460
rect 279187 477395 279253 477396
rect 278451 477052 278517 477053
rect 278451 476988 278452 477052
rect 278516 476988 278517 477052
rect 278451 476987 278517 476988
rect 280846 476237 280906 479710
rect 283422 476237 283482 479710
rect 285998 477053 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293358 479710 293508 479770
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 285995 477052 286061 477053
rect 285995 476988 285996 477052
rect 286060 476988 286061 477052
rect 285995 476987 286061 476988
rect 288206 476781 288266 479710
rect 288203 476780 288269 476781
rect 288203 476716 288204 476780
rect 288268 476716 288269 476780
rect 288203 476715 288269 476716
rect 290966 476509 291026 479710
rect 290963 476508 291029 476509
rect 290963 476444 290964 476508
rect 291028 476444 291029 476508
rect 290963 476443 291029 476444
rect 293358 476237 293418 479710
rect 295934 476237 295994 479710
rect 298510 476373 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 305960 479710 306114 479770
rect 308544 479710 308690 479770
rect 310992 479710 311082 479770
rect 300902 476781 300962 479710
rect 300899 476780 300965 476781
rect 300899 476716 300900 476780
rect 300964 476716 300965 476780
rect 300899 476715 300965 476716
rect 303478 476373 303538 479710
rect 306054 476509 306114 479710
rect 308630 476645 308690 479710
rect 311022 477189 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318472 479770 318532 480080
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 318472 479710 318626 479770
rect 320920 479710 321018 479770
rect 311019 477188 311085 477189
rect 311019 477124 311020 477188
rect 311084 477124 311085 477188
rect 311019 477123 311085 477124
rect 313414 476645 313474 479710
rect 315806 476781 315866 479710
rect 318566 476781 318626 479710
rect 320958 476917 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 323350 477053 323410 479710
rect 325926 477053 325986 479710
rect 323347 477052 323413 477053
rect 323347 476988 323348 477052
rect 323412 476988 323413 477052
rect 323347 476987 323413 476988
rect 325923 477052 325989 477053
rect 325923 476988 325924 477052
rect 325988 476988 325989 477052
rect 325923 476987 325989 476988
rect 320955 476916 321021 476917
rect 320955 476852 320956 476916
rect 321020 476852 321021 476916
rect 320955 476851 321021 476852
rect 315803 476780 315869 476781
rect 315803 476716 315804 476780
rect 315868 476716 315869 476780
rect 315803 476715 315869 476716
rect 318563 476780 318629 476781
rect 318563 476716 318564 476780
rect 318628 476716 318629 476780
rect 318563 476715 318629 476716
rect 308627 476644 308693 476645
rect 308627 476580 308628 476644
rect 308692 476580 308693 476644
rect 308627 476579 308693 476580
rect 313411 476644 313477 476645
rect 313411 476580 313412 476644
rect 313476 476580 313477 476644
rect 313411 476579 313477 476580
rect 306051 476508 306117 476509
rect 306051 476444 306052 476508
rect 306116 476444 306117 476508
rect 306051 476443 306117 476444
rect 298507 476372 298573 476373
rect 298507 476308 298508 476372
rect 298572 476308 298573 476372
rect 298507 476307 298573 476308
rect 303475 476372 303541 476373
rect 303475 476308 303476 476372
rect 303540 476308 303541 476372
rect 303475 476307 303541 476308
rect 248275 476236 248341 476237
rect 248275 476172 248276 476236
rect 248340 476172 248341 476236
rect 248275 476171 248341 476172
rect 250667 476236 250733 476237
rect 250667 476172 250668 476236
rect 250732 476172 250733 476236
rect 250667 476171 250733 476172
rect 253611 476236 253677 476237
rect 253611 476172 253612 476236
rect 253676 476172 253677 476236
rect 253611 476171 253677 476172
rect 258395 476236 258461 476237
rect 258395 476172 258396 476236
rect 258460 476172 258461 476236
rect 258395 476171 258461 476172
rect 260971 476236 261037 476237
rect 260971 476172 260972 476236
rect 261036 476172 261037 476236
rect 260971 476171 261037 476172
rect 263547 476236 263613 476237
rect 263547 476172 263548 476236
rect 263612 476172 263613 476236
rect 263547 476171 263613 476172
rect 265939 476236 266005 476237
rect 265939 476172 265940 476236
rect 266004 476172 266005 476236
rect 265939 476171 266005 476172
rect 268331 476236 268397 476237
rect 268331 476172 268332 476236
rect 268396 476172 268397 476236
rect 268331 476171 268397 476172
rect 273483 476236 273549 476237
rect 273483 476172 273484 476236
rect 273548 476172 273549 476236
rect 273483 476171 273549 476172
rect 276059 476236 276125 476237
rect 276059 476172 276060 476236
rect 276124 476172 276125 476236
rect 276059 476171 276125 476172
rect 280843 476236 280909 476237
rect 280843 476172 280844 476236
rect 280908 476172 280909 476236
rect 280843 476171 280909 476172
rect 283419 476236 283485 476237
rect 283419 476172 283420 476236
rect 283484 476172 283485 476236
rect 283419 476171 283485 476172
rect 293355 476236 293421 476237
rect 293355 476172 293356 476236
rect 293420 476172 293421 476236
rect 293355 476171 293421 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 350947 445772 351013 445773
rect 350947 445708 350948 445772
rect 351012 445708 351013 445772
rect 350947 445707 351013 445708
rect 350950 443730 351010 445707
rect 350840 443670 351010 443730
rect 350840 443202 350900 443670
rect 220272 439174 220620 439206
rect 220272 438938 220328 439174
rect 220564 438938 220620 439174
rect 220272 438854 220620 438938
rect 220272 438618 220328 438854
rect 220564 438618 220620 438854
rect 220272 438586 220620 438618
rect 356000 439174 356348 439206
rect 356000 438938 356056 439174
rect 356292 438938 356348 439174
rect 356000 438854 356348 438938
rect 356000 438618 356056 438854
rect 356292 438618 356348 438854
rect 356000 438586 356348 438618
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 403174 220620 403206
rect 220272 402938 220328 403174
rect 220564 402938 220620 403174
rect 220272 402854 220620 402938
rect 220272 402618 220328 402854
rect 220564 402618 220620 402854
rect 220272 402586 220620 402618
rect 356000 403174 356348 403206
rect 356000 402938 356056 403174
rect 356292 402938 356348 403174
rect 356000 402854 356348 402938
rect 356000 402618 356056 402854
rect 356292 402618 356348 402854
rect 356000 402586 356348 402618
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 220272 367174 220620 367206
rect 220272 366938 220328 367174
rect 220564 366938 220620 367174
rect 220272 366854 220620 366938
rect 220272 366618 220328 366854
rect 220564 366618 220620 366854
rect 220272 366586 220620 366618
rect 356000 367174 356348 367206
rect 356000 366938 356056 367174
rect 356292 366938 356348 367174
rect 356000 366854 356348 366938
rect 356000 366618 356056 366854
rect 356292 366618 356348 366854
rect 356000 366586 356348 366618
rect 220952 363454 221300 363486
rect 220952 363218 221008 363454
rect 221244 363218 221300 363454
rect 220952 363134 221300 363218
rect 220952 362898 221008 363134
rect 221244 362898 221300 363134
rect 220952 362866 221300 362898
rect 355320 363454 355668 363486
rect 355320 363218 355376 363454
rect 355612 363218 355668 363454
rect 355320 363134 355668 363218
rect 355320 362898 355376 363134
rect 355612 362898 355668 363134
rect 355320 362866 355668 362898
rect 236056 359410 236116 360060
rect 235950 359350 236116 359410
rect 237144 359410 237204 360060
rect 238232 359410 238292 360060
rect 239592 359818 239652 360060
rect 238894 359758 239652 359818
rect 240544 359818 240604 360060
rect 241768 359818 241828 360060
rect 243128 359818 243188 360060
rect 240544 359758 240978 359818
rect 241768 359758 241898 359818
rect 238894 359410 238954 359758
rect 237144 359350 237298 359410
rect 238232 359350 238402 359410
rect 235950 358597 236010 359350
rect 235947 358596 236013 358597
rect 235947 358532 235948 358596
rect 236012 358532 236013 358596
rect 235947 358531 236013 358532
rect 221514 331174 222134 358064
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 219939 289100 220005 289101
rect 219939 289036 219940 289100
rect 220004 289036 220005 289100
rect 219939 289035 220005 289036
rect 218651 282844 218717 282845
rect 218651 282780 218652 282844
rect 218716 282780 218717 282844
rect 218651 282779 218717 282780
rect 219755 282844 219821 282845
rect 219755 282780 219756 282844
rect 219820 282780 219821 282844
rect 219755 282779 219821 282780
rect 221514 281537 222134 294618
rect 225234 334894 225854 358064
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 281537 225854 298338
rect 228954 338614 229574 358064
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 281537 229574 302058
rect 232674 342334 233294 358064
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232674 306334 233294 341778
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232674 281537 233294 305778
rect 236394 346054 237014 358064
rect 237238 356285 237298 359350
rect 238342 357237 238402 359350
rect 238526 359350 238954 359410
rect 238526 357370 238586 359350
rect 238526 357310 238954 357370
rect 238339 357236 238405 357237
rect 238339 357172 238340 357236
rect 238404 357172 238405 357236
rect 238339 357171 238405 357172
rect 238894 357101 238954 357310
rect 238891 357100 238957 357101
rect 238891 357036 238892 357100
rect 238956 357036 238957 357100
rect 238891 357035 238957 357036
rect 237235 356284 237301 356285
rect 237235 356220 237236 356284
rect 237300 356220 237301 356284
rect 237235 356219 237301 356220
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 236394 310054 237014 345498
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 236394 281537 237014 309498
rect 240114 349774 240734 357940
rect 240918 356149 240978 359758
rect 241838 356829 241898 359758
rect 243126 359758 243188 359818
rect 244216 359818 244276 360060
rect 245440 359818 245500 360060
rect 246528 359818 246588 360060
rect 247616 359818 247676 360060
rect 248296 359818 248356 360060
rect 248704 359818 248764 360060
rect 244216 359758 244658 359818
rect 245440 359758 245578 359818
rect 246528 359758 246682 359818
rect 243126 357373 243186 359758
rect 243123 357372 243189 357373
rect 243123 357308 243124 357372
rect 243188 357308 243189 357372
rect 243123 357307 243189 357308
rect 241835 356828 241901 356829
rect 241835 356764 241836 356828
rect 241900 356764 241901 356828
rect 241835 356763 241901 356764
rect 240915 356148 240981 356149
rect 240915 356084 240916 356148
rect 240980 356084 240981 356148
rect 240915 356083 240981 356084
rect 240114 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 240734 349774
rect 240114 349454 240734 349538
rect 240114 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 240734 349454
rect 240114 313774 240734 349218
rect 240114 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 240734 313774
rect 240114 313454 240734 313538
rect 240114 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 240734 313454
rect 240114 281537 240734 313218
rect 243834 353494 244454 357940
rect 244598 356965 244658 359758
rect 244595 356964 244661 356965
rect 244595 356900 244596 356964
rect 244660 356900 244661 356964
rect 244595 356899 244661 356900
rect 245518 356693 245578 359758
rect 245515 356692 245581 356693
rect 245515 356628 245516 356692
rect 245580 356628 245581 356692
rect 245515 356627 245581 356628
rect 246622 356421 246682 359758
rect 247542 359758 247676 359818
rect 248278 359758 248356 359818
rect 248646 359758 248764 359818
rect 250064 359818 250124 360060
rect 250744 359818 250804 360060
rect 251288 359818 251348 360060
rect 252376 359818 252436 360060
rect 253464 359818 253524 360060
rect 250064 359758 250178 359818
rect 247542 356557 247602 359758
rect 248278 357373 248338 359758
rect 248646 357373 248706 359758
rect 248275 357372 248341 357373
rect 248275 357308 248276 357372
rect 248340 357308 248341 357372
rect 248275 357307 248341 357308
rect 248643 357372 248709 357373
rect 248643 357308 248644 357372
rect 248708 357308 248709 357372
rect 248643 357307 248709 357308
rect 250118 356693 250178 359758
rect 250670 359758 250804 359818
rect 251222 359758 251348 359818
rect 252326 359758 252436 359818
rect 253430 359758 253524 359818
rect 253600 359818 253660 360060
rect 254552 359818 254612 360060
rect 255912 359818 255972 360060
rect 253600 359758 253674 359818
rect 250670 357373 250730 359758
rect 251222 357373 251282 359758
rect 250667 357372 250733 357373
rect 250667 357308 250668 357372
rect 250732 357308 250733 357372
rect 250667 357307 250733 357308
rect 251219 357372 251285 357373
rect 251219 357308 251220 357372
rect 251284 357308 251285 357372
rect 251219 357307 251285 357308
rect 252326 356693 252386 359758
rect 250115 356692 250181 356693
rect 250115 356628 250116 356692
rect 250180 356628 250181 356692
rect 250115 356627 250181 356628
rect 252323 356692 252389 356693
rect 252323 356628 252324 356692
rect 252388 356628 252389 356692
rect 252323 356627 252389 356628
rect 253430 356557 253490 359758
rect 253614 357373 253674 359758
rect 254534 359758 254612 359818
rect 255822 359758 255972 359818
rect 253611 357372 253677 357373
rect 253611 357308 253612 357372
rect 253676 357308 253677 357372
rect 253611 357307 253677 357308
rect 247539 356556 247605 356557
rect 247539 356492 247540 356556
rect 247604 356492 247605 356556
rect 247539 356491 247605 356492
rect 253427 356556 253493 356557
rect 253427 356492 253428 356556
rect 253492 356492 253493 356556
rect 253427 356491 253493 356492
rect 246619 356420 246685 356421
rect 246619 356356 246620 356420
rect 246684 356356 246685 356420
rect 246619 356355 246685 356356
rect 243834 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 244454 353494
rect 243834 353174 244454 353258
rect 243834 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 244454 353174
rect 243834 317494 244454 352938
rect 243834 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 244454 317494
rect 243834 317174 244454 317258
rect 243834 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 244454 317174
rect 243834 281537 244454 316938
rect 253794 327454 254414 358064
rect 254534 357373 254594 359758
rect 254531 357372 254597 357373
rect 254531 357308 254532 357372
rect 254596 357308 254597 357372
rect 254531 357307 254597 357308
rect 255822 356693 255882 359758
rect 256048 359410 256108 360060
rect 257000 359818 257060 360060
rect 257000 359758 257170 359818
rect 256006 359350 256108 359410
rect 256006 357373 256066 359350
rect 257110 357373 257170 359758
rect 258088 359410 258148 360060
rect 258496 359410 258556 360060
rect 258088 359350 258274 359410
rect 256003 357372 256069 357373
rect 256003 357308 256004 357372
rect 256068 357308 256069 357372
rect 256003 357307 256069 357308
rect 257107 357372 257173 357373
rect 257107 357308 257108 357372
rect 257172 357308 257173 357372
rect 257107 357307 257173 357308
rect 255819 356692 255885 356693
rect 255819 356628 255820 356692
rect 255884 356628 255885 356692
rect 255819 356627 255885 356628
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 281537 254414 290898
rect 257514 331174 258134 357940
rect 258214 356690 258274 359350
rect 258398 359350 258556 359410
rect 259448 359410 259508 360060
rect 260672 359410 260732 360060
rect 261080 359410 261140 360060
rect 259448 359350 259562 359410
rect 258398 357373 258458 359350
rect 258395 357372 258461 357373
rect 258395 357308 258396 357372
rect 258460 357308 258461 357372
rect 258395 357307 258461 357308
rect 259502 356693 259562 359350
rect 260606 359350 260732 359410
rect 260974 359350 261140 359410
rect 261760 359410 261820 360060
rect 262848 359410 262908 360060
rect 261760 359350 262138 359410
rect 258395 356692 258461 356693
rect 258395 356690 258396 356692
rect 258214 356630 258396 356690
rect 258395 356628 258396 356630
rect 258460 356628 258461 356692
rect 258395 356627 258461 356628
rect 259499 356692 259565 356693
rect 259499 356628 259500 356692
rect 259564 356628 259565 356692
rect 259499 356627 259565 356628
rect 260606 356421 260666 359350
rect 260974 357373 261034 359350
rect 260971 357372 261037 357373
rect 260971 357308 260972 357372
rect 261036 357308 261037 357372
rect 260971 357307 261037 357308
rect 260603 356420 260669 356421
rect 260603 356356 260604 356420
rect 260668 356356 260669 356420
rect 260603 356355 260669 356356
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 281537 258134 294618
rect 261234 334894 261854 357940
rect 262078 357373 262138 359350
rect 262814 359350 262908 359410
rect 263528 359410 263588 360060
rect 263936 359410 263996 360060
rect 263528 359350 263610 359410
rect 262814 357373 262874 359350
rect 263550 357373 263610 359350
rect 263918 359350 263996 359410
rect 265296 359410 265356 360060
rect 265976 359410 266036 360060
rect 266384 359410 266444 360060
rect 267608 359410 267668 360060
rect 268288 359546 268348 360060
rect 268696 359546 268756 360060
rect 268288 359486 268394 359546
rect 265296 359350 265818 359410
rect 263918 357373 263978 359350
rect 262075 357372 262141 357373
rect 262075 357308 262076 357372
rect 262140 357308 262141 357372
rect 262075 357307 262141 357308
rect 262811 357372 262877 357373
rect 262811 357308 262812 357372
rect 262876 357308 262877 357372
rect 262811 357307 262877 357308
rect 263547 357372 263613 357373
rect 263547 357308 263548 357372
rect 263612 357308 263613 357372
rect 263547 357307 263613 357308
rect 263915 357372 263981 357373
rect 263915 357308 263916 357372
rect 263980 357308 263981 357372
rect 263915 357307 263981 357308
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 281537 261854 298338
rect 264954 338614 265574 357940
rect 265758 357373 265818 359350
rect 265942 359350 266036 359410
rect 266310 359350 266444 359410
rect 267598 359350 267668 359410
rect 265755 357372 265821 357373
rect 265755 357308 265756 357372
rect 265820 357308 265821 357372
rect 265755 357307 265821 357308
rect 265942 356557 266002 359350
rect 266310 357373 266370 359350
rect 267598 357373 267658 359350
rect 268334 357373 268394 359486
rect 268518 359486 268756 359546
rect 269784 359546 269844 360060
rect 271008 359546 271068 360060
rect 269784 359486 269866 359546
rect 268518 357373 268578 359486
rect 266307 357372 266373 357373
rect 266307 357308 266308 357372
rect 266372 357308 266373 357372
rect 266307 357307 266373 357308
rect 267595 357372 267661 357373
rect 267595 357308 267596 357372
rect 267660 357308 267661 357372
rect 267595 357307 267661 357308
rect 268331 357372 268397 357373
rect 268331 357308 268332 357372
rect 268396 357308 268397 357372
rect 268331 357307 268397 357308
rect 268515 357372 268581 357373
rect 268515 357308 268516 357372
rect 268580 357308 268581 357372
rect 268515 357307 268581 357308
rect 265939 356556 266005 356557
rect 265939 356492 265940 356556
rect 266004 356492 266005 356556
rect 265939 356491 266005 356492
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 281537 265574 302058
rect 268674 342334 269294 357940
rect 269806 357373 269866 359486
rect 270910 359486 271068 359546
rect 270910 357373 270970 359486
rect 271144 359410 271204 360060
rect 272232 359546 272292 360060
rect 271094 359350 271204 359410
rect 272198 359486 272292 359546
rect 271094 357373 271154 359350
rect 272198 357373 272258 359486
rect 273320 359410 273380 360060
rect 273592 359410 273652 360060
rect 274408 359410 274468 360060
rect 273302 359350 273380 359410
rect 273486 359350 273652 359410
rect 274406 359350 274468 359410
rect 275768 359410 275828 360060
rect 276040 359410 276100 360060
rect 276992 359410 277052 360060
rect 275768 359350 275938 359410
rect 276040 359350 276122 359410
rect 269803 357372 269869 357373
rect 269803 357308 269804 357372
rect 269868 357308 269869 357372
rect 269803 357307 269869 357308
rect 270907 357372 270973 357373
rect 270907 357308 270908 357372
rect 270972 357308 270973 357372
rect 270907 357307 270973 357308
rect 271091 357372 271157 357373
rect 271091 357308 271092 357372
rect 271156 357308 271157 357372
rect 271091 357307 271157 357308
rect 272195 357372 272261 357373
rect 272195 357308 272196 357372
rect 272260 357308 272261 357372
rect 272195 357307 272261 357308
rect 268674 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 269294 342334
rect 268674 342014 269294 342098
rect 268674 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 269294 342014
rect 268674 306334 269294 341778
rect 268674 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 269294 306334
rect 268674 306014 269294 306098
rect 268674 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 269294 306014
rect 268674 281537 269294 305778
rect 272394 346054 273014 358064
rect 273302 357373 273362 359350
rect 273299 357372 273365 357373
rect 273299 357308 273300 357372
rect 273364 357308 273365 357372
rect 273299 357307 273365 357308
rect 273486 356149 273546 359350
rect 274406 357373 274466 359350
rect 275878 357373 275938 359350
rect 276062 358189 276122 359350
rect 276982 359350 277052 359410
rect 278080 359410 278140 360060
rect 278488 359410 278548 360060
rect 278080 359350 278146 359410
rect 276059 358188 276125 358189
rect 276059 358124 276060 358188
rect 276124 358124 276125 358188
rect 276059 358123 276125 358124
rect 274403 357372 274469 357373
rect 274403 357308 274404 357372
rect 274468 357308 274469 357372
rect 274403 357307 274469 357308
rect 275875 357372 275941 357373
rect 275875 357308 275876 357372
rect 275940 357308 275941 357372
rect 275875 357307 275941 357308
rect 273483 356148 273549 356149
rect 273483 356084 273484 356148
rect 273548 356084 273549 356148
rect 273483 356083 273549 356084
rect 272394 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 273014 346054
rect 272394 345734 273014 345818
rect 272394 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 273014 345734
rect 272394 310054 273014 345498
rect 272394 309818 272426 310054
rect 272662 309818 272746 310054
rect 272982 309818 273014 310054
rect 272394 309734 273014 309818
rect 272394 309498 272426 309734
rect 272662 309498 272746 309734
rect 272982 309498 273014 309734
rect 272394 281537 273014 309498
rect 276114 349774 276734 357940
rect 276982 357373 277042 359350
rect 276979 357372 277045 357373
rect 276979 357308 276980 357372
rect 277044 357308 277045 357372
rect 276979 357307 277045 357308
rect 278086 356693 278146 359350
rect 278454 359350 278548 359410
rect 279168 359410 279228 360060
rect 280936 359410 280996 360060
rect 283520 359546 283580 360060
rect 279168 359350 279250 359410
rect 278083 356692 278149 356693
rect 278083 356628 278084 356692
rect 278148 356628 278149 356692
rect 278083 356627 278149 356628
rect 278454 356149 278514 359350
rect 279190 356557 279250 359350
rect 280846 359350 280996 359410
rect 283422 359486 283580 359546
rect 285968 359546 286028 360060
rect 285968 359486 286058 359546
rect 279187 356556 279253 356557
rect 279187 356492 279188 356556
rect 279252 356492 279253 356556
rect 279187 356491 279253 356492
rect 278451 356148 278517 356149
rect 278451 356084 278452 356148
rect 278516 356084 278517 356148
rect 278451 356083 278517 356084
rect 276114 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 276734 349774
rect 276114 349454 276734 349538
rect 276114 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 276734 349454
rect 276114 313774 276734 349218
rect 276114 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 276734 313774
rect 276114 313454 276734 313538
rect 276114 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 276734 313454
rect 276114 281537 276734 313218
rect 279834 353494 280454 358064
rect 280846 356149 280906 359350
rect 283422 357373 283482 359486
rect 285998 357373 286058 359486
rect 288280 359410 288340 360060
rect 291000 359410 291060 360060
rect 293448 359410 293508 360060
rect 288206 359350 288340 359410
rect 290966 359350 291060 359410
rect 293358 359350 293508 359410
rect 295896 359410 295956 360060
rect 298480 359410 298540 360060
rect 300928 359410 300988 360060
rect 303512 359410 303572 360060
rect 305960 359410 306020 360060
rect 308544 359410 308604 360060
rect 295896 359350 295994 359410
rect 298480 359350 298570 359410
rect 288206 357373 288266 359350
rect 283419 357372 283485 357373
rect 283419 357308 283420 357372
rect 283484 357308 283485 357372
rect 283419 357307 283485 357308
rect 285995 357372 286061 357373
rect 285995 357308 285996 357372
rect 286060 357308 286061 357372
rect 285995 357307 286061 357308
rect 288203 357372 288269 357373
rect 288203 357308 288204 357372
rect 288268 357308 288269 357372
rect 288203 357307 288269 357308
rect 280843 356148 280909 356149
rect 280843 356084 280844 356148
rect 280908 356084 280909 356148
rect 280843 356083 280909 356084
rect 279834 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 280454 353494
rect 279834 353174 280454 353258
rect 279834 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 280454 353174
rect 279834 317494 280454 352938
rect 279834 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 280454 317494
rect 279834 317174 280454 317258
rect 279834 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 280454 317174
rect 279834 281537 280454 316938
rect 289794 327454 290414 358064
rect 290966 357373 291026 359350
rect 293358 357373 293418 359350
rect 290963 357372 291029 357373
rect 290963 357308 290964 357372
rect 291028 357308 291029 357372
rect 290963 357307 291029 357308
rect 293355 357372 293421 357373
rect 293355 357308 293356 357372
rect 293420 357308 293421 357372
rect 293355 357307 293421 357308
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 281537 290414 290898
rect 293514 331174 294134 357940
rect 295934 357373 295994 359350
rect 295931 357372 295997 357373
rect 295931 357308 295932 357372
rect 295996 357308 295997 357372
rect 295931 357307 295997 357308
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 281537 294134 294618
rect 297234 334894 297854 358064
rect 298510 357373 298570 359350
rect 300902 359350 300988 359410
rect 303478 359350 303572 359410
rect 305870 359350 306020 359410
rect 308078 359350 308604 359410
rect 310992 359410 311052 360060
rect 313440 359410 313500 360060
rect 315888 359410 315948 360060
rect 318472 359410 318532 360060
rect 310992 359350 311082 359410
rect 300902 358189 300962 359350
rect 300899 358188 300965 358189
rect 300899 358124 300900 358188
rect 300964 358124 300965 358188
rect 300899 358123 300965 358124
rect 298507 357372 298573 357373
rect 298507 357308 298508 357372
rect 298572 357308 298573 357372
rect 298507 357307 298573 357308
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 201008 259174 201328 259206
rect 201008 258938 201050 259174
rect 201286 258938 201328 259174
rect 201008 258854 201328 258938
rect 201008 258618 201050 258854
rect 201286 258618 201328 258854
rect 201008 258586 201328 258618
rect 231728 259174 232048 259206
rect 231728 258938 231770 259174
rect 232006 258938 232048 259174
rect 231728 258854 232048 258938
rect 231728 258618 231770 258854
rect 232006 258618 232048 258854
rect 231728 258586 232048 258618
rect 262448 259174 262768 259206
rect 262448 258938 262490 259174
rect 262726 258938 262768 259174
rect 262448 258854 262768 258938
rect 262448 258618 262490 258854
rect 262726 258618 262768 258854
rect 262448 258586 262768 258618
rect 293168 259174 293488 259206
rect 293168 258938 293210 259174
rect 293446 258938 293488 259174
rect 293168 258854 293488 258938
rect 293168 258618 293210 258854
rect 293446 258618 293488 258854
rect 293168 258586 293488 258618
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 216368 255454 216688 255486
rect 216368 255218 216410 255454
rect 216646 255218 216688 255454
rect 216368 255134 216688 255218
rect 216368 254898 216410 255134
rect 216646 254898 216688 255134
rect 216368 254866 216688 254898
rect 247088 255454 247408 255486
rect 247088 255218 247130 255454
rect 247366 255218 247408 255454
rect 247088 255134 247408 255218
rect 247088 254898 247130 255134
rect 247366 254898 247408 255134
rect 247088 254866 247408 254898
rect 277808 255454 278128 255486
rect 277808 255218 277850 255454
rect 278086 255218 278128 255454
rect 277808 255134 278128 255218
rect 277808 254898 277850 255134
rect 278086 254898 278128 255134
rect 277808 254866 278128 254898
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 201008 223174 201328 223206
rect 201008 222938 201050 223174
rect 201286 222938 201328 223174
rect 201008 222854 201328 222938
rect 201008 222618 201050 222854
rect 201286 222618 201328 222854
rect 201008 222586 201328 222618
rect 231728 223174 232048 223206
rect 231728 222938 231770 223174
rect 232006 222938 232048 223174
rect 231728 222854 232048 222938
rect 231728 222618 231770 222854
rect 232006 222618 232048 222854
rect 231728 222586 232048 222618
rect 262448 223174 262768 223206
rect 262448 222938 262490 223174
rect 262726 222938 262768 223174
rect 262448 222854 262768 222938
rect 262448 222618 262490 222854
rect 262726 222618 262768 222854
rect 262448 222586 262768 222618
rect 293168 223174 293488 223206
rect 293168 222938 293210 223174
rect 293446 222938 293488 223174
rect 293168 222854 293488 222938
rect 293168 222618 293210 222854
rect 293446 222618 293488 222854
rect 293168 222586 293488 222618
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 216368 219454 216688 219486
rect 216368 219218 216410 219454
rect 216646 219218 216688 219454
rect 216368 219134 216688 219218
rect 216368 218898 216410 219134
rect 216646 218898 216688 219134
rect 216368 218866 216688 218898
rect 247088 219454 247408 219486
rect 247088 219218 247130 219454
rect 247366 219218 247408 219454
rect 247088 219134 247408 219218
rect 247088 218898 247130 219134
rect 247366 218898 247408 219134
rect 247088 218866 247408 218898
rect 277808 219454 278128 219486
rect 277808 219218 277850 219454
rect 278086 219218 278128 219454
rect 277808 219134 278128 219218
rect 277808 218898 277850 219134
rect 278086 218898 278128 219134
rect 277808 218866 278128 218898
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 201008 187174 201328 187206
rect 201008 186938 201050 187174
rect 201286 186938 201328 187174
rect 201008 186854 201328 186938
rect 201008 186618 201050 186854
rect 201286 186618 201328 186854
rect 201008 186586 201328 186618
rect 231728 187174 232048 187206
rect 231728 186938 231770 187174
rect 232006 186938 232048 187174
rect 231728 186854 232048 186938
rect 231728 186618 231770 186854
rect 232006 186618 232048 186854
rect 231728 186586 232048 186618
rect 262448 187174 262768 187206
rect 262448 186938 262490 187174
rect 262726 186938 262768 187174
rect 262448 186854 262768 186938
rect 262448 186618 262490 186854
rect 262726 186618 262768 186854
rect 262448 186586 262768 186618
rect 293168 187174 293488 187206
rect 293168 186938 293210 187174
rect 293446 186938 293488 187174
rect 293168 186854 293488 186938
rect 293168 186618 293210 186854
rect 293446 186618 293488 186854
rect 293168 186586 293488 186618
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 185648 183454 185968 183486
rect 185648 183218 185690 183454
rect 185926 183218 185968 183454
rect 185648 183134 185968 183218
rect 185648 182898 185690 183134
rect 185926 182898 185968 183134
rect 185648 182866 185968 182898
rect 216368 183454 216688 183486
rect 216368 183218 216410 183454
rect 216646 183218 216688 183454
rect 216368 183134 216688 183218
rect 216368 182898 216410 183134
rect 216646 182898 216688 183134
rect 216368 182866 216688 182898
rect 247088 183454 247408 183486
rect 247088 183218 247130 183454
rect 247366 183218 247408 183454
rect 247088 183134 247408 183218
rect 247088 182898 247130 183134
rect 247366 182898 247408 183134
rect 247088 182866 247408 182898
rect 277808 183454 278128 183486
rect 277808 183218 277850 183454
rect 278086 183218 278128 183454
rect 277808 183134 278128 183218
rect 277808 182898 277850 183134
rect 278086 182898 278128 183134
rect 277808 182866 278128 182898
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 201008 151174 201328 151206
rect 201008 150938 201050 151174
rect 201286 150938 201328 151174
rect 201008 150854 201328 150938
rect 201008 150618 201050 150854
rect 201286 150618 201328 150854
rect 201008 150586 201328 150618
rect 231728 151174 232048 151206
rect 231728 150938 231770 151174
rect 232006 150938 232048 151174
rect 231728 150854 232048 150938
rect 231728 150618 231770 150854
rect 232006 150618 232048 150854
rect 231728 150586 232048 150618
rect 262448 151174 262768 151206
rect 262448 150938 262490 151174
rect 262726 150938 262768 151174
rect 262448 150854 262768 150938
rect 262448 150618 262490 150854
rect 262726 150618 262768 150854
rect 262448 150586 262768 150618
rect 293168 151174 293488 151206
rect 293168 150938 293210 151174
rect 293446 150938 293488 151174
rect 293168 150854 293488 150938
rect 293168 150618 293210 150854
rect 293446 150618 293488 150854
rect 293168 150586 293488 150618
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 185648 147454 185968 147486
rect 185648 147218 185690 147454
rect 185926 147218 185968 147454
rect 185648 147134 185968 147218
rect 185648 146898 185690 147134
rect 185926 146898 185968 147134
rect 185648 146866 185968 146898
rect 216368 147454 216688 147486
rect 216368 147218 216410 147454
rect 216646 147218 216688 147454
rect 216368 147134 216688 147218
rect 216368 146898 216410 147134
rect 216646 146898 216688 147134
rect 216368 146866 216688 146898
rect 247088 147454 247408 147486
rect 247088 147218 247130 147454
rect 247366 147218 247408 147454
rect 247088 147134 247408 147218
rect 247088 146898 247130 147134
rect 247366 146898 247408 147134
rect 247088 146866 247408 146898
rect 277808 147454 278128 147486
rect 277808 147218 277850 147454
rect 278086 147218 278128 147454
rect 277808 147134 278128 147218
rect 277808 146898 277850 147134
rect 278086 146898 278128 147134
rect 277808 146866 278128 146898
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 201008 115174 201328 115206
rect 201008 114938 201050 115174
rect 201286 114938 201328 115174
rect 201008 114854 201328 114938
rect 201008 114618 201050 114854
rect 201286 114618 201328 114854
rect 201008 114586 201328 114618
rect 231728 115174 232048 115206
rect 231728 114938 231770 115174
rect 232006 114938 232048 115174
rect 231728 114854 232048 114938
rect 231728 114618 231770 114854
rect 232006 114618 232048 114854
rect 231728 114586 232048 114618
rect 262448 115174 262768 115206
rect 262448 114938 262490 115174
rect 262726 114938 262768 115174
rect 262448 114854 262768 114938
rect 262448 114618 262490 114854
rect 262726 114618 262768 114854
rect 262448 114586 262768 114618
rect 293168 115174 293488 115206
rect 293168 114938 293210 115174
rect 293446 114938 293488 115174
rect 293168 114854 293488 114938
rect 293168 114618 293210 114854
rect 293446 114618 293488 114854
rect 293168 114586 293488 114618
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 216368 111454 216688 111486
rect 216368 111218 216410 111454
rect 216646 111218 216688 111454
rect 216368 111134 216688 111218
rect 216368 110898 216410 111134
rect 216646 110898 216688 111134
rect 216368 110866 216688 110898
rect 247088 111454 247408 111486
rect 247088 111218 247130 111454
rect 247366 111218 247408 111454
rect 247088 111134 247408 111218
rect 247088 110898 247130 111134
rect 247366 110898 247408 111134
rect 247088 110866 247408 110898
rect 277808 111454 278128 111486
rect 277808 111218 277850 111454
rect 278086 111218 278128 111454
rect 277808 111134 278128 111218
rect 277808 110898 277850 111134
rect 278086 110898 278128 111134
rect 277808 110866 278128 110898
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 79174 186134 79743
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 79743
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 50614 193574 79743
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 54334 197294 79743
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 58054 201014 79743
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 61774 204734 79743
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 65494 208454 79743
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 75454 218414 79743
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 79174 222134 79743
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 79743
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 50614 229574 79743
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 54334 233294 79743
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 58054 237014 79743
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 61774 240734 79743
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 65494 244454 79743
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 75454 254414 79743
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 79174 258134 79743
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 79743
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 50614 265574 79743
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 54334 269294 79743
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 58054 273014 79743
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 61774 276734 79743
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 276114 25774 276734 61218
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 65494 280454 79743
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 279834 29494 280454 64938
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 75454 290414 79743
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 79174 294134 79743
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 338614 301574 357940
rect 303478 357373 303538 359350
rect 303475 357372 303541 357373
rect 303475 357308 303476 357372
rect 303540 357308 303541 357372
rect 303475 357307 303541 357308
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 342334 305294 358064
rect 305870 357373 305930 359350
rect 308078 357373 308138 359350
rect 305867 357372 305933 357373
rect 305867 357308 305868 357372
rect 305932 357308 305933 357372
rect 305867 357307 305933 357308
rect 308075 357372 308141 357373
rect 308075 357308 308076 357372
rect 308140 357308 308141 357372
rect 308075 357307 308141 357308
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 304674 306334 305294 341778
rect 304674 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 305294 306334
rect 304674 306014 305294 306098
rect 304674 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 305294 306014
rect 304674 270334 305294 305778
rect 308394 346054 309014 357940
rect 311022 357373 311082 359350
rect 313414 359350 313500 359410
rect 315622 359350 315948 359410
rect 318382 359350 318532 359410
rect 320920 359410 320980 360060
rect 323368 359410 323428 360060
rect 325952 359410 326012 360060
rect 320920 359350 321018 359410
rect 311019 357372 311085 357373
rect 311019 357308 311020 357372
rect 311084 357308 311085 357372
rect 311019 357307 311085 357308
rect 308394 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 309014 346054
rect 308394 345734 309014 345818
rect 308394 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 309014 345734
rect 308394 310054 309014 345498
rect 308394 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 309014 310054
rect 308394 309734 309014 309818
rect 308394 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 309014 309734
rect 308394 279580 309014 309498
rect 312114 349774 312734 358064
rect 313414 357373 313474 359350
rect 315622 357373 315682 359350
rect 313411 357372 313477 357373
rect 313411 357308 313412 357372
rect 313476 357308 313477 357372
rect 313411 357307 313477 357308
rect 315619 357372 315685 357373
rect 315619 357308 315620 357372
rect 315684 357308 315685 357372
rect 315619 357307 315685 357308
rect 312114 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 312734 349774
rect 312114 349454 312734 349538
rect 312114 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 312734 349454
rect 312114 313774 312734 349218
rect 312114 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 312734 313774
rect 312114 313454 312734 313538
rect 312114 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 312734 313454
rect 304674 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 305294 270334
rect 304674 270014 305294 270098
rect 304674 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 305294 270014
rect 304674 234334 305294 269778
rect 312114 277774 312734 313218
rect 312114 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 312734 277774
rect 312114 277454 312734 277538
rect 312114 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 312734 277454
rect 308528 255454 308848 255486
rect 308528 255218 308570 255454
rect 308806 255218 308848 255454
rect 308528 255134 308848 255218
rect 308528 254898 308570 255134
rect 308806 254898 308848 255134
rect 308528 254866 308848 254898
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 304674 198334 305294 233778
rect 312114 241774 312734 277218
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 308528 219454 308848 219486
rect 308528 219218 308570 219454
rect 308806 219218 308848 219454
rect 308528 219134 308848 219218
rect 308528 218898 308570 219134
rect 308806 218898 308848 219134
rect 308528 218866 308848 218898
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 304674 162334 305294 197778
rect 312114 205774 312734 241218
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 308528 183454 308848 183486
rect 308528 183218 308570 183454
rect 308806 183218 308848 183454
rect 308528 183134 308848 183218
rect 308528 182898 308570 183134
rect 308806 182898 308848 183134
rect 308528 182866 308848 182898
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 312114 169774 312734 205218
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 308528 147454 308848 147486
rect 308528 147218 308570 147454
rect 308806 147218 308848 147454
rect 308528 147134 308848 147218
rect 308528 146898 308570 147134
rect 308806 146898 308848 147134
rect 308528 146866 308848 146898
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304674 90334 305294 125778
rect 312114 133774 312734 169218
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 308528 111454 308848 111486
rect 308528 111218 308570 111454
rect 308806 111218 308848 111454
rect 308528 111134 308848 111218
rect 308528 110898 308570 111134
rect 308806 110898 308848 111134
rect 308528 110866 308848 110898
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 304674 54334 305294 89778
rect 312114 97774 312734 133218
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 58054 309014 80068
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 61774 312734 97218
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 312114 25774 312734 61218
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 353494 316454 357940
rect 318382 357373 318442 359350
rect 320958 357373 321018 359350
rect 323350 359350 323428 359410
rect 325926 359350 326012 359410
rect 318379 357372 318445 357373
rect 318379 357308 318380 357372
rect 318444 357308 318445 357372
rect 318379 357307 318445 357308
rect 320955 357372 321021 357373
rect 320955 357308 320956 357372
rect 321020 357308 321021 357372
rect 320955 357307 321021 357308
rect 323350 356149 323410 359350
rect 325926 358733 325986 359350
rect 325923 358732 325989 358733
rect 325923 358668 325924 358732
rect 325988 358668 325989 358732
rect 325923 358667 325989 358668
rect 323347 356148 323413 356149
rect 323347 356084 323348 356148
rect 323412 356084 323413 356148
rect 323347 356083 323413 356084
rect 315834 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 316454 353494
rect 315834 353174 316454 353258
rect 315834 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 316454 353174
rect 315834 317494 316454 352938
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 315834 281494 316454 316938
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 315834 245494 316454 280938
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 101494 316454 136938
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 315834 65494 316454 100938
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 327454 326414 357940
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 331174 330134 358064
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 334894 333854 358064
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 338614 337574 358064
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 342334 341294 358064
rect 340674 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 341294 342334
rect 340674 342014 341294 342098
rect 340674 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 341294 342014
rect 340674 306334 341294 341778
rect 340674 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 341294 306334
rect 340674 306014 341294 306098
rect 340674 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 341294 306014
rect 340674 270334 341294 305778
rect 340674 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 341294 270334
rect 340674 270014 341294 270098
rect 340674 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 341294 270014
rect 340674 234334 341294 269778
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 340674 162334 341294 197778
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 340674 126334 341294 161778
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 90334 341294 125778
rect 340674 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 341294 90334
rect 340674 90014 341294 90098
rect 340674 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 341294 90014
rect 340674 54334 341294 89778
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 346054 345014 358064
rect 344394 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 345014 346054
rect 344394 345734 345014 345818
rect 344394 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 345014 345734
rect 344394 310054 345014 345498
rect 344394 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 345014 310054
rect 344394 309734 345014 309818
rect 344394 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 345014 309734
rect 344394 274054 345014 309498
rect 344394 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 345014 274054
rect 344394 273734 345014 273818
rect 344394 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 345014 273734
rect 344394 238054 345014 273498
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 344394 166054 345014 201498
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 344394 130054 345014 165498
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 344394 94054 345014 129498
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 344394 58054 345014 93498
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 349774 348734 358064
rect 348114 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 348734 349774
rect 348114 349454 348734 349538
rect 348114 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 348734 349454
rect 348114 313774 348734 349218
rect 348114 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 348734 313774
rect 348114 313454 348734 313538
rect 348114 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 348734 313454
rect 348114 277774 348734 313218
rect 348114 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 348734 277774
rect 348114 277454 348734 277538
rect 348114 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 348734 277454
rect 348114 241774 348734 277218
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 97774 348734 133218
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 353494 352454 358064
rect 351834 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 352454 353494
rect 351834 353174 352454 353258
rect 351834 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 352454 353174
rect 351834 317494 352454 352938
rect 351834 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 352454 317494
rect 351834 317174 352454 317258
rect 351834 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 352454 317174
rect 351834 281494 352454 316938
rect 356654 297397 356714 596939
rect 357022 298757 357082 597075
rect 357574 359549 357634 597347
rect 357571 359548 357637 359549
rect 357571 359484 357572 359548
rect 357636 359484 357637 359548
rect 357571 359483 357637 359484
rect 357019 298756 357085 298757
rect 357019 298692 357020 298756
rect 357084 298692 357085 298756
rect 357019 298691 357085 298692
rect 356651 297396 356717 297397
rect 356651 297332 356652 297396
rect 356716 297332 356717 297396
rect 356651 297331 356717 297332
rect 357942 294541 358002 607411
rect 358859 597276 358925 597277
rect 358859 597212 358860 597276
rect 358924 597212 358925 597276
rect 358859 597211 358925 597212
rect 358123 592652 358189 592653
rect 358123 592588 358124 592652
rect 358188 592588 358189 592652
rect 358123 592587 358189 592588
rect 357939 294540 358005 294541
rect 357939 294476 357940 294540
rect 358004 294476 358005 294540
rect 357939 294475 358005 294476
rect 358126 282301 358186 592587
rect 358862 359413 358922 597211
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 359411 487252 359477 487253
rect 359411 487188 359412 487252
rect 359476 487188 359477 487252
rect 359411 487187 359477 487188
rect 358859 359412 358925 359413
rect 358859 359348 358860 359412
rect 358924 359348 358925 359412
rect 358859 359347 358925 359348
rect 359414 293181 359474 487187
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 359411 293180 359477 293181
rect 359411 293116 359412 293180
rect 359476 293116 359477 293180
rect 359411 293115 359477 293116
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 358123 282300 358189 282301
rect 358123 282236 358124 282300
rect 358188 282236 358189 282300
rect 358123 282235 358189 282236
rect 351834 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 352454 281494
rect 351834 281174 352454 281258
rect 351834 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 352454 281174
rect 351834 245494 352454 280938
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351834 101494 352454 136938
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 364208 219454 364528 219486
rect 364208 219218 364250 219454
rect 364486 219218 364528 219454
rect 364208 219134 364528 219218
rect 364208 218898 364250 219134
rect 364486 218898 364528 219134
rect 364208 218866 364528 218898
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 364208 183454 364528 183486
rect 364208 183218 364250 183454
rect 364486 183218 364528 183454
rect 364208 183134 364528 183218
rect 364208 182898 364250 183134
rect 364486 182898 364528 183134
rect 364208 182866 364528 182898
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 364208 147454 364528 147486
rect 364208 147218 364250 147454
rect 364486 147218 364528 147454
rect 364208 147134 364528 147218
rect 364208 146898 364250 147134
rect 364486 146898 364528 147134
rect 364208 146866 364528 146898
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 364208 111454 364528 111486
rect 364208 111218 364250 111454
rect 364486 111218 364528 111454
rect 364208 111134 364528 111218
rect 364208 110898 364250 111134
rect 364486 110898 364528 111134
rect 364208 110866 364528 110898
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 364208 75454 364528 75486
rect 364208 75218 364250 75454
rect 364486 75218 364528 75454
rect 364208 75134 364528 75218
rect 364208 74898 364250 75134
rect 364486 74898 364528 75134
rect 364208 74866 364528 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 379568 223174 379888 223206
rect 379568 222938 379610 223174
rect 379846 222938 379888 223174
rect 379568 222854 379888 222938
rect 379568 222618 379610 222854
rect 379846 222618 379888 222854
rect 379568 222586 379888 222618
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 379568 187174 379888 187206
rect 379568 186938 379610 187174
rect 379846 186938 379888 187174
rect 379568 186854 379888 186938
rect 379568 186618 379610 186854
rect 379846 186618 379888 186854
rect 379568 186586 379888 186618
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 379568 151174 379888 151206
rect 379568 150938 379610 151174
rect 379846 150938 379888 151174
rect 379568 150854 379888 150938
rect 379568 150618 379610 150854
rect 379846 150618 379888 150854
rect 379568 150586 379888 150618
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 379568 115174 379888 115206
rect 379568 114938 379610 115174
rect 379846 114938 379888 115174
rect 379568 114854 379888 114938
rect 379568 114618 379610 114854
rect 379846 114618 379888 114854
rect 379568 114586 379888 114618
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 379568 79174 379888 79206
rect 379568 78938 379610 79174
rect 379846 78938 379888 79174
rect 379568 78854 379888 78938
rect 379568 78618 379610 78854
rect 379846 78618 379888 78854
rect 379568 78586 379888 78618
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 395291 700500 395357 700501
rect 395291 700436 395292 700500
rect 395356 700436 395357 700500
rect 395291 700435 395357 700436
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 395294 351117 395354 700435
rect 397499 699820 397565 699821
rect 397499 699756 397500 699820
rect 397564 699756 397565 699820
rect 397499 699755 397565 699756
rect 397131 513772 397197 513773
rect 397131 513708 397132 513772
rect 397196 513708 397197 513772
rect 397131 513707 397197 513708
rect 397134 394637 397194 513707
rect 397315 487388 397381 487389
rect 397315 487324 397316 487388
rect 397380 487324 397381 487388
rect 397315 487323 397381 487324
rect 397318 446453 397378 487323
rect 397315 446452 397381 446453
rect 397315 446388 397316 446452
rect 397380 446388 397381 446452
rect 397315 446387 397381 446388
rect 397131 394636 397197 394637
rect 397131 394572 397132 394636
rect 397196 394572 397197 394636
rect 397131 394571 397197 394572
rect 397318 368389 397378 446387
rect 397315 368388 397381 368389
rect 397315 368324 397316 368388
rect 397380 368324 397381 368388
rect 397315 368323 397381 368324
rect 397502 352613 397562 699755
rect 397794 687454 398414 704282
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 398603 700364 398669 700365
rect 398603 700300 398604 700364
rect 398668 700300 398669 700364
rect 398603 700299 398669 700300
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 685244 398414 686898
rect 397499 352612 397565 352613
rect 397499 352548 397500 352612
rect 397564 352548 397565 352612
rect 397499 352547 397565 352548
rect 395291 351116 395357 351117
rect 395291 351052 395292 351116
rect 395356 351052 395357 351116
rect 395291 351051 395357 351052
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 397794 327454 398414 358064
rect 398606 349757 398666 700299
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 685244 402134 690618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 685244 405854 694338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 685244 409574 698058
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 685244 434414 686898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 685244 438134 690618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 685244 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 685244 445574 698058
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 685244 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 685244 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 685244 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 685244 481574 698058
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 685244 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 685244 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 685244 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 685244 517574 698058
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 530899 685948 530965 685949
rect 530899 685884 530900 685948
rect 530964 685884 530965 685948
rect 530899 685883 530965 685884
rect 530902 683770 530962 685883
rect 530840 683710 530962 683770
rect 530840 683202 530900 683710
rect 400272 655174 400620 655206
rect 400272 654938 400328 655174
rect 400564 654938 400620 655174
rect 400272 654854 400620 654938
rect 400272 654618 400328 654854
rect 400564 654618 400620 654854
rect 400272 654586 400620 654618
rect 536000 655174 536348 655206
rect 536000 654938 536056 655174
rect 536292 654938 536348 655174
rect 536000 654854 536348 654938
rect 536000 654618 536056 654854
rect 536292 654618 536348 654854
rect 536000 654586 536348 654618
rect 400952 651454 401300 651486
rect 400952 651218 401008 651454
rect 401244 651218 401300 651454
rect 400952 651134 401300 651218
rect 400952 650898 401008 651134
rect 401244 650898 401300 651134
rect 400952 650866 401300 650898
rect 535320 651454 535668 651486
rect 535320 651218 535376 651454
rect 535612 651218 535668 651454
rect 535320 651134 535668 651218
rect 535320 650898 535376 651134
rect 535612 650898 535668 651134
rect 535320 650866 535668 650898
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 400272 619174 400620 619206
rect 400272 618938 400328 619174
rect 400564 618938 400620 619174
rect 400272 618854 400620 618938
rect 400272 618618 400328 618854
rect 400564 618618 400620 618854
rect 400272 618586 400620 618618
rect 536000 619174 536348 619206
rect 536000 618938 536056 619174
rect 536292 618938 536348 619174
rect 536000 618854 536348 618938
rect 536000 618618 536056 618854
rect 536292 618618 536348 618854
rect 536000 618586 536348 618618
rect 400952 615454 401300 615486
rect 400952 615218 401008 615454
rect 401244 615218 401300 615454
rect 400952 615134 401300 615218
rect 400952 614898 401008 615134
rect 401244 614898 401300 615134
rect 400952 614866 401300 614898
rect 535320 615454 535668 615486
rect 535320 615218 535376 615454
rect 535612 615218 535668 615454
rect 535320 615134 535668 615218
rect 535320 614898 535376 615134
rect 535612 614898 535668 615134
rect 535320 614866 535668 614898
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 416056 599450 416116 600100
rect 417144 599450 417204 600100
rect 418232 599450 418292 600100
rect 419592 599450 419652 600100
rect 420544 599450 420604 600100
rect 416056 599390 416146 599450
rect 417144 599390 417250 599450
rect 418232 599390 418354 599450
rect 416086 597549 416146 599390
rect 417190 597549 417250 599390
rect 418294 597549 418354 599390
rect 419582 599390 419652 599450
rect 420502 599390 420604 599450
rect 421768 599450 421828 600100
rect 423128 599450 423188 600100
rect 424216 599450 424276 600100
rect 421768 599390 421850 599450
rect 416083 597548 416149 597549
rect 416083 597484 416084 597548
rect 416148 597484 416149 597548
rect 416083 597483 416149 597484
rect 417187 597548 417253 597549
rect 417187 597484 417188 597548
rect 417252 597484 417253 597548
rect 417187 597483 417253 597484
rect 418291 597548 418357 597549
rect 418291 597484 418292 597548
rect 418356 597484 418357 597548
rect 418291 597483 418357 597484
rect 419582 596733 419642 599390
rect 420502 597549 420562 599390
rect 421790 597549 421850 599390
rect 423078 599390 423188 599450
rect 424182 599390 424276 599450
rect 425440 599450 425500 600100
rect 426528 599450 426588 600100
rect 427616 599450 427676 600100
rect 428296 599450 428356 600100
rect 428704 599450 428764 600100
rect 425440 599390 425530 599450
rect 426528 599390 426634 599450
rect 427616 599390 427738 599450
rect 423078 597549 423138 599390
rect 424182 597549 424242 599390
rect 425470 597549 425530 599390
rect 426574 597549 426634 599390
rect 427678 597549 427738 599390
rect 428230 599390 428356 599450
rect 428598 599390 428764 599450
rect 430064 599450 430124 600100
rect 430744 599450 430804 600100
rect 431288 599450 431348 600100
rect 432376 599450 432436 600100
rect 433464 599450 433524 600100
rect 430064 599390 430130 599450
rect 420499 597548 420565 597549
rect 420499 597484 420500 597548
rect 420564 597484 420565 597548
rect 420499 597483 420565 597484
rect 421787 597548 421853 597549
rect 421787 597484 421788 597548
rect 421852 597484 421853 597548
rect 421787 597483 421853 597484
rect 423075 597548 423141 597549
rect 423075 597484 423076 597548
rect 423140 597484 423141 597548
rect 423075 597483 423141 597484
rect 424179 597548 424245 597549
rect 424179 597484 424180 597548
rect 424244 597484 424245 597548
rect 424179 597483 424245 597484
rect 425467 597548 425533 597549
rect 425467 597484 425468 597548
rect 425532 597484 425533 597548
rect 425467 597483 425533 597484
rect 426571 597548 426637 597549
rect 426571 597484 426572 597548
rect 426636 597484 426637 597548
rect 426571 597483 426637 597484
rect 427675 597548 427741 597549
rect 427675 597484 427676 597548
rect 427740 597484 427741 597548
rect 427675 597483 427741 597484
rect 428230 596733 428290 599390
rect 428598 597549 428658 599390
rect 430070 597549 430130 599390
rect 430622 599390 430804 599450
rect 431174 599390 431348 599450
rect 431726 599390 432436 599450
rect 433382 599390 433524 599450
rect 433600 599450 433660 600100
rect 434552 599450 434612 600100
rect 435912 599589 435972 600100
rect 435909 599588 435975 599589
rect 435909 599524 435910 599588
rect 435974 599524 435975 599588
rect 435909 599523 435975 599524
rect 436048 599450 436108 600100
rect 433600 599390 433810 599450
rect 430622 597549 430682 599390
rect 428595 597548 428661 597549
rect 428595 597484 428596 597548
rect 428660 597484 428661 597548
rect 428595 597483 428661 597484
rect 430067 597548 430133 597549
rect 430067 597484 430068 597548
rect 430132 597484 430133 597548
rect 430067 597483 430133 597484
rect 430619 597548 430685 597549
rect 430619 597484 430620 597548
rect 430684 597484 430685 597548
rect 430619 597483 430685 597484
rect 431174 596733 431234 599390
rect 419579 596732 419645 596733
rect 419579 596668 419580 596732
rect 419644 596668 419645 596732
rect 419579 596667 419645 596668
rect 428227 596732 428293 596733
rect 428227 596668 428228 596732
rect 428292 596668 428293 596732
rect 428227 596667 428293 596668
rect 431171 596732 431237 596733
rect 431171 596668 431172 596732
rect 431236 596668 431237 596732
rect 431726 596730 431786 599390
rect 433382 596733 433442 599390
rect 433750 597549 433810 599390
rect 434486 599390 434612 599450
rect 435958 599390 436108 599450
rect 437000 599450 437060 600100
rect 438088 599450 438148 600100
rect 437000 599390 437122 599450
rect 434486 597549 434546 599390
rect 435958 597549 436018 599390
rect 437062 597549 437122 599390
rect 437982 599390 438148 599450
rect 438496 599450 438556 600100
rect 439448 599450 439508 600100
rect 440672 599450 440732 600100
rect 441080 599450 441140 600100
rect 441760 599450 441820 600100
rect 442848 599450 442908 600100
rect 443528 599450 443588 600100
rect 443936 599450 443996 600100
rect 438496 599390 438594 599450
rect 439448 599390 439514 599450
rect 440672 599390 440802 599450
rect 441080 599390 441170 599450
rect 437982 597549 438042 599390
rect 433747 597548 433813 597549
rect 433747 597484 433748 597548
rect 433812 597484 433813 597548
rect 433747 597483 433813 597484
rect 434483 597548 434549 597549
rect 434483 597484 434484 597548
rect 434548 597484 434549 597548
rect 434483 597483 434549 597484
rect 435955 597548 436021 597549
rect 435955 597484 435956 597548
rect 436020 597484 436021 597548
rect 435955 597483 436021 597484
rect 437059 597548 437125 597549
rect 437059 597484 437060 597548
rect 437124 597484 437125 597548
rect 437059 597483 437125 597484
rect 437979 597548 438045 597549
rect 437979 597484 437980 597548
rect 438044 597484 438045 597548
rect 437979 597483 438045 597484
rect 438534 597141 438594 599390
rect 439454 597549 439514 599390
rect 439451 597548 439517 597549
rect 439451 597484 439452 597548
rect 439516 597484 439517 597548
rect 439451 597483 439517 597484
rect 440742 597141 440802 599390
rect 438531 597140 438597 597141
rect 438531 597076 438532 597140
rect 438596 597076 438597 597140
rect 438531 597075 438597 597076
rect 440739 597140 440805 597141
rect 440739 597076 440740 597140
rect 440804 597076 440805 597140
rect 440739 597075 440805 597076
rect 441110 597005 441170 599390
rect 441662 599390 441820 599450
rect 442766 599390 442908 599450
rect 443502 599390 443588 599450
rect 443870 599390 443996 599450
rect 445296 599450 445356 600100
rect 445976 599450 446036 600100
rect 446384 599450 446444 600100
rect 447608 599450 447668 600100
rect 448288 599450 448348 600100
rect 448696 599450 448756 600100
rect 449784 599450 449844 600100
rect 450859 599588 450925 599589
rect 450859 599524 450860 599588
rect 450924 599524 450925 599588
rect 450859 599523 450925 599524
rect 445296 599390 445402 599450
rect 441662 597005 441722 599390
rect 442766 597549 442826 599390
rect 443502 597549 443562 599390
rect 443870 597549 443930 599390
rect 445342 597549 445402 599390
rect 445894 599390 446036 599450
rect 446262 599390 446444 599450
rect 447550 599390 447668 599450
rect 448286 599390 448348 599450
rect 448654 599390 448756 599450
rect 449758 599390 449844 599450
rect 445894 597549 445954 599390
rect 442763 597548 442829 597549
rect 442763 597484 442764 597548
rect 442828 597484 442829 597548
rect 442763 597483 442829 597484
rect 443499 597548 443565 597549
rect 443499 597484 443500 597548
rect 443564 597484 443565 597548
rect 443499 597483 443565 597484
rect 443867 597548 443933 597549
rect 443867 597484 443868 597548
rect 443932 597484 443933 597548
rect 443867 597483 443933 597484
rect 445339 597548 445405 597549
rect 445339 597484 445340 597548
rect 445404 597484 445405 597548
rect 445339 597483 445405 597484
rect 445891 597548 445957 597549
rect 445891 597484 445892 597548
rect 445956 597484 445957 597548
rect 445891 597483 445957 597484
rect 446262 597005 446322 599390
rect 447550 597005 447610 599390
rect 448286 597549 448346 599390
rect 448283 597548 448349 597549
rect 448283 597484 448284 597548
rect 448348 597484 448349 597548
rect 448283 597483 448349 597484
rect 448654 597005 448714 599390
rect 441107 597004 441173 597005
rect 441107 596940 441108 597004
rect 441172 596940 441173 597004
rect 441107 596939 441173 596940
rect 441659 597004 441725 597005
rect 441659 596940 441660 597004
rect 441724 596940 441725 597004
rect 441659 596939 441725 596940
rect 446259 597004 446325 597005
rect 446259 596940 446260 597004
rect 446324 596940 446325 597004
rect 446259 596939 446325 596940
rect 447547 597004 447613 597005
rect 447547 596940 447548 597004
rect 447612 596940 447613 597004
rect 447547 596939 447613 596940
rect 448651 597004 448717 597005
rect 448651 596940 448652 597004
rect 448716 596940 448717 597004
rect 448651 596939 448717 596940
rect 431907 596732 431973 596733
rect 431907 596730 431908 596732
rect 431726 596670 431908 596730
rect 431171 596667 431237 596668
rect 431907 596668 431908 596670
rect 431972 596668 431973 596732
rect 431907 596667 431973 596668
rect 433379 596732 433445 596733
rect 433379 596668 433380 596732
rect 433444 596668 433445 596732
rect 433379 596667 433445 596668
rect 449758 596325 449818 599390
rect 450862 596461 450922 599523
rect 451008 599450 451068 600100
rect 451144 599589 451204 600100
rect 451141 599588 451207 599589
rect 451141 599524 451142 599588
rect 451206 599524 451207 599588
rect 452232 599586 452292 600100
rect 453320 599586 453380 600100
rect 451141 599523 451207 599524
rect 452150 599526 452292 599586
rect 453254 599526 453380 599586
rect 453592 599586 453652 600100
rect 454408 599586 454468 600100
rect 455768 599586 455828 600100
rect 456040 599586 456100 600100
rect 456992 599586 457052 600100
rect 458080 599586 458140 600100
rect 458488 599586 458548 600100
rect 459168 599586 459228 600100
rect 453592 599526 453682 599586
rect 452150 599453 452210 599526
rect 452147 599452 452213 599453
rect 451008 599390 451106 599450
rect 451046 597549 451106 599390
rect 452147 599388 452148 599452
rect 452212 599388 452213 599452
rect 452147 599387 452213 599388
rect 451043 597548 451109 597549
rect 451043 597484 451044 597548
rect 451108 597484 451109 597548
rect 451043 597483 451109 597484
rect 453254 597413 453314 599526
rect 453251 597412 453317 597413
rect 453251 597348 453252 597412
rect 453316 597348 453317 597412
rect 453251 597347 453317 597348
rect 453622 596597 453682 599526
rect 454358 599526 454468 599586
rect 455646 599526 455828 599586
rect 456014 599526 456100 599586
rect 456934 599526 457052 599586
rect 458038 599526 458140 599586
rect 458406 599526 458548 599586
rect 459142 599526 459228 599586
rect 454358 597005 454418 599526
rect 455646 597005 455706 599526
rect 456014 597549 456074 599526
rect 456011 597548 456077 597549
rect 456011 597484 456012 597548
rect 456076 597484 456077 597548
rect 456011 597483 456077 597484
rect 454355 597004 454421 597005
rect 454355 596940 454356 597004
rect 454420 596940 454421 597004
rect 454355 596939 454421 596940
rect 455643 597004 455709 597005
rect 455643 596940 455644 597004
rect 455708 596940 455709 597004
rect 455643 596939 455709 596940
rect 453619 596596 453685 596597
rect 453619 596532 453620 596596
rect 453684 596532 453685 596596
rect 453619 596531 453685 596532
rect 450859 596460 450925 596461
rect 450859 596396 450860 596460
rect 450924 596396 450925 596460
rect 450859 596395 450925 596396
rect 456934 596325 456994 599526
rect 458038 596733 458098 599526
rect 458406 596869 458466 599526
rect 459142 597141 459202 599526
rect 460936 599450 460996 600100
rect 463520 599450 463580 600100
rect 465968 599450 466028 600100
rect 468280 599450 468340 600100
rect 471000 599450 471060 600100
rect 460936 599390 461042 599450
rect 463520 599390 463618 599450
rect 460982 597277 461042 599390
rect 463558 597549 463618 599390
rect 465950 599390 466028 599450
rect 468158 599390 468340 599450
rect 470366 599390 471060 599450
rect 473448 599450 473508 600100
rect 475896 599450 475956 600100
rect 478480 599450 478540 600100
rect 480928 599450 480988 600100
rect 483512 599450 483572 600100
rect 473448 599390 473554 599450
rect 465950 597549 466010 599390
rect 468158 597549 468218 599390
rect 463555 597548 463621 597549
rect 463555 597484 463556 597548
rect 463620 597484 463621 597548
rect 463555 597483 463621 597484
rect 465947 597548 466013 597549
rect 465947 597484 465948 597548
rect 466012 597484 466013 597548
rect 465947 597483 466013 597484
rect 468155 597548 468221 597549
rect 468155 597484 468156 597548
rect 468220 597484 468221 597548
rect 468155 597483 468221 597484
rect 460979 597276 461045 597277
rect 460979 597212 460980 597276
rect 461044 597212 461045 597276
rect 460979 597211 461045 597212
rect 459139 597140 459205 597141
rect 459139 597076 459140 597140
rect 459204 597076 459205 597140
rect 459139 597075 459205 597076
rect 458403 596868 458469 596869
rect 458403 596804 458404 596868
rect 458468 596804 458469 596868
rect 458403 596803 458469 596804
rect 458035 596732 458101 596733
rect 458035 596668 458036 596732
rect 458100 596668 458101 596732
rect 458035 596667 458101 596668
rect 470366 596325 470426 599390
rect 473494 597549 473554 599390
rect 475886 599390 475956 599450
rect 478462 599390 478540 599450
rect 480854 599390 480988 599450
rect 483430 599390 483572 599450
rect 485960 599450 486020 600100
rect 488544 599450 488604 600100
rect 490992 599450 491052 600100
rect 493440 599450 493500 600100
rect 485960 599390 486066 599450
rect 488544 599390 488642 599450
rect 475886 597549 475946 599390
rect 478462 597549 478522 599390
rect 473491 597548 473557 597549
rect 473491 597484 473492 597548
rect 473556 597484 473557 597548
rect 473491 597483 473557 597484
rect 475883 597548 475949 597549
rect 475883 597484 475884 597548
rect 475948 597484 475949 597548
rect 475883 597483 475949 597484
rect 478459 597548 478525 597549
rect 478459 597484 478460 597548
rect 478524 597484 478525 597548
rect 478459 597483 478525 597484
rect 480854 597005 480914 599390
rect 483430 597549 483490 599390
rect 486006 597549 486066 599390
rect 488582 597549 488642 599390
rect 489686 599390 491052 599450
rect 493366 599390 493500 599450
rect 495888 599450 495948 600100
rect 498472 599450 498532 600100
rect 500920 599450 500980 600100
rect 503368 599450 503428 600100
rect 505952 599450 506012 600100
rect 495888 599390 496002 599450
rect 498472 599390 498578 599450
rect 483427 597548 483493 597549
rect 483427 597484 483428 597548
rect 483492 597484 483493 597548
rect 483427 597483 483493 597484
rect 486003 597548 486069 597549
rect 486003 597484 486004 597548
rect 486068 597484 486069 597548
rect 486003 597483 486069 597484
rect 488579 597548 488645 597549
rect 488579 597484 488580 597548
rect 488644 597484 488645 597548
rect 488579 597483 488645 597484
rect 480851 597004 480917 597005
rect 480851 596940 480852 597004
rect 480916 596940 480917 597004
rect 480851 596939 480917 596940
rect 489686 596325 489746 599390
rect 493366 596733 493426 599390
rect 495942 597549 496002 599390
rect 498518 597549 498578 599390
rect 500910 599390 500980 599450
rect 503302 599390 503428 599450
rect 505878 599390 506012 599450
rect 500910 597549 500970 599390
rect 495939 597548 496005 597549
rect 495939 597484 495940 597548
rect 496004 597484 496005 597548
rect 495939 597483 496005 597484
rect 498515 597548 498581 597549
rect 498515 597484 498516 597548
rect 498580 597484 498581 597548
rect 498515 597483 498581 597484
rect 500907 597548 500973 597549
rect 500907 597484 500908 597548
rect 500972 597484 500973 597548
rect 500907 597483 500973 597484
rect 503302 597005 503362 599390
rect 503299 597004 503365 597005
rect 503299 596940 503300 597004
rect 503364 596940 503365 597004
rect 503299 596939 503365 596940
rect 505878 596869 505938 599390
rect 505875 596868 505941 596869
rect 505875 596804 505876 596868
rect 505940 596804 505941 596868
rect 505875 596803 505941 596804
rect 493363 596732 493429 596733
rect 493363 596668 493364 596732
rect 493428 596668 493429 596732
rect 493363 596667 493429 596668
rect 449755 596324 449821 596325
rect 449755 596260 449756 596324
rect 449820 596260 449821 596324
rect 449755 596259 449821 596260
rect 456931 596324 456997 596325
rect 456931 596260 456932 596324
rect 456996 596260 456997 596324
rect 456931 596259 456997 596260
rect 470363 596324 470429 596325
rect 470363 596260 470364 596324
rect 470428 596260 470429 596324
rect 470363 596259 470429 596260
rect 489683 596324 489749 596325
rect 489683 596260 489684 596324
rect 489748 596260 489749 596324
rect 489683 596259 489749 596260
rect 399339 594556 399405 594557
rect 399339 594492 399340 594556
rect 399404 594492 399405 594556
rect 399339 594491 399405 594492
rect 398787 444276 398853 444277
rect 398787 444212 398788 444276
rect 398852 444212 398853 444276
rect 398787 444211 398853 444212
rect 398603 349756 398669 349757
rect 398603 349692 398604 349756
rect 398668 349692 398669 349756
rect 398603 349691 398669 349692
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 398790 311133 398850 444211
rect 399342 348397 399402 594491
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 530899 565860 530965 565861
rect 530899 565796 530900 565860
rect 530964 565796 530965 565860
rect 530899 565795 530965 565796
rect 530902 564090 530962 565795
rect 530840 564030 530962 564090
rect 530840 563202 530900 564030
rect 400272 547174 400620 547206
rect 400272 546938 400328 547174
rect 400564 546938 400620 547174
rect 400272 546854 400620 546938
rect 400272 546618 400328 546854
rect 400564 546618 400620 546854
rect 400272 546586 400620 546618
rect 536000 547174 536348 547206
rect 536000 546938 536056 547174
rect 536292 546938 536348 547174
rect 536000 546854 536348 546938
rect 536000 546618 536056 546854
rect 536292 546618 536348 546854
rect 536000 546586 536348 546618
rect 400952 543454 401300 543486
rect 400952 543218 401008 543454
rect 401244 543218 401300 543454
rect 400952 543134 401300 543218
rect 400952 542898 401008 543134
rect 401244 542898 401300 543134
rect 400952 542866 401300 542898
rect 535320 543454 535668 543486
rect 535320 543218 535376 543454
rect 535612 543218 535668 543454
rect 535320 543134 535668 543218
rect 535320 542898 535376 543134
rect 535612 542898 535668 543134
rect 535320 542866 535668 542898
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 400272 511174 400620 511206
rect 400272 510938 400328 511174
rect 400564 510938 400620 511174
rect 400272 510854 400620 510938
rect 400272 510618 400328 510854
rect 400564 510618 400620 510854
rect 400272 510586 400620 510618
rect 536000 511174 536348 511206
rect 536000 510938 536056 511174
rect 536292 510938 536348 511174
rect 536000 510854 536348 510938
rect 536000 510618 536056 510854
rect 536292 510618 536348 510854
rect 536000 510586 536348 510618
rect 400952 507454 401300 507486
rect 400952 507218 401008 507454
rect 401244 507218 401300 507454
rect 400952 507134 401300 507218
rect 400952 506898 401008 507134
rect 401244 506898 401300 507134
rect 400952 506866 401300 506898
rect 535320 507454 535668 507486
rect 535320 507218 535376 507454
rect 535612 507218 535668 507454
rect 535320 507134 535668 507218
rect 535320 506898 535376 507134
rect 535612 506898 535668 507134
rect 535320 506866 535668 506898
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 416056 479770 416116 480080
rect 417144 479770 417204 480080
rect 418232 479770 418292 480080
rect 419592 479770 419652 480080
rect 420544 479770 420604 480080
rect 416056 479710 416146 479770
rect 417144 479710 417250 479770
rect 418232 479710 418354 479770
rect 416086 477461 416146 479710
rect 417190 477461 417250 479710
rect 418294 477461 418354 479710
rect 419582 479710 419652 479770
rect 420502 479710 420604 479770
rect 421768 479770 421828 480080
rect 423128 479770 423188 480080
rect 424216 479770 424276 480080
rect 421768 479710 421850 479770
rect 416083 477460 416149 477461
rect 416083 477396 416084 477460
rect 416148 477396 416149 477460
rect 416083 477395 416149 477396
rect 417187 477460 417253 477461
rect 417187 477396 417188 477460
rect 417252 477396 417253 477460
rect 417187 477395 417253 477396
rect 418291 477460 418357 477461
rect 418291 477396 418292 477460
rect 418356 477396 418357 477460
rect 418291 477395 418357 477396
rect 419582 476509 419642 479710
rect 420502 477461 420562 479710
rect 421790 477461 421850 479710
rect 423078 479710 423188 479770
rect 424182 479710 424276 479770
rect 425440 479770 425500 480080
rect 426528 479770 426588 480080
rect 427616 479770 427676 480080
rect 428296 479770 428356 480080
rect 428704 479770 428764 480080
rect 425440 479710 425530 479770
rect 426528 479710 426634 479770
rect 427616 479710 427738 479770
rect 423078 477461 423138 479710
rect 424182 477461 424242 479710
rect 425470 477461 425530 479710
rect 426574 477461 426634 479710
rect 427678 477461 427738 479710
rect 428230 479710 428356 479770
rect 428598 479710 428764 479770
rect 430064 479770 430124 480080
rect 430744 479770 430804 480080
rect 430064 479710 430130 479770
rect 420499 477460 420565 477461
rect 420499 477396 420500 477460
rect 420564 477396 420565 477460
rect 420499 477395 420565 477396
rect 421787 477460 421853 477461
rect 421787 477396 421788 477460
rect 421852 477396 421853 477460
rect 421787 477395 421853 477396
rect 423075 477460 423141 477461
rect 423075 477396 423076 477460
rect 423140 477396 423141 477460
rect 423075 477395 423141 477396
rect 424179 477460 424245 477461
rect 424179 477396 424180 477460
rect 424244 477396 424245 477460
rect 424179 477395 424245 477396
rect 425467 477460 425533 477461
rect 425467 477396 425468 477460
rect 425532 477396 425533 477460
rect 425467 477395 425533 477396
rect 426571 477460 426637 477461
rect 426571 477396 426572 477460
rect 426636 477396 426637 477460
rect 426571 477395 426637 477396
rect 427675 477460 427741 477461
rect 427675 477396 427676 477460
rect 427740 477396 427741 477460
rect 427675 477395 427741 477396
rect 419579 476508 419645 476509
rect 419579 476444 419580 476508
rect 419644 476444 419645 476508
rect 419579 476443 419645 476444
rect 428230 476237 428290 479710
rect 428598 478413 428658 479710
rect 430070 478413 430130 479710
rect 430622 479710 430804 479770
rect 431288 479770 431348 480080
rect 432376 479770 432436 480080
rect 433464 479770 433524 480080
rect 431288 479710 431418 479770
rect 432376 479710 432522 479770
rect 428595 478412 428661 478413
rect 428595 478348 428596 478412
rect 428660 478348 428661 478412
rect 428595 478347 428661 478348
rect 430067 478412 430133 478413
rect 430067 478348 430068 478412
rect 430132 478348 430133 478412
rect 430067 478347 430133 478348
rect 430622 476237 430682 479710
rect 431358 478277 431418 479710
rect 432462 478277 432522 479710
rect 433382 479710 433524 479770
rect 433600 479770 433660 480080
rect 434552 479770 434612 480080
rect 435912 479770 435972 480080
rect 433600 479710 433810 479770
rect 431355 478276 431421 478277
rect 431355 478212 431356 478276
rect 431420 478212 431421 478276
rect 431355 478211 431421 478212
rect 432459 478276 432525 478277
rect 432459 478212 432460 478276
rect 432524 478212 432525 478276
rect 432459 478211 432525 478212
rect 433382 477461 433442 479710
rect 433379 477460 433445 477461
rect 433379 477396 433380 477460
rect 433444 477396 433445 477460
rect 433379 477395 433445 477396
rect 433750 476509 433810 479710
rect 434486 479710 434612 479770
rect 435774 479710 435972 479770
rect 434486 477461 434546 479710
rect 435774 477461 435834 479710
rect 436048 479090 436108 480080
rect 437000 479770 437060 480080
rect 438088 479770 438148 480080
rect 438496 479770 438556 480080
rect 439448 479770 439508 480080
rect 440672 479770 440732 480080
rect 441080 479770 441140 480080
rect 441760 479770 441820 480080
rect 442848 479770 442908 480080
rect 443528 479770 443588 480080
rect 443936 479770 443996 480080
rect 437000 479710 437122 479770
rect 438088 479710 438226 479770
rect 438496 479710 438594 479770
rect 439448 479710 439514 479770
rect 440672 479710 440802 479770
rect 441080 479710 441170 479770
rect 435958 479030 436108 479090
rect 434483 477460 434549 477461
rect 434483 477396 434484 477460
rect 434548 477396 434549 477460
rect 434483 477395 434549 477396
rect 435771 477460 435837 477461
rect 435771 477396 435772 477460
rect 435836 477396 435837 477460
rect 435771 477395 435837 477396
rect 435958 477189 436018 479030
rect 437062 477461 437122 479710
rect 438166 477461 438226 479710
rect 437059 477460 437125 477461
rect 437059 477396 437060 477460
rect 437124 477396 437125 477460
rect 437059 477395 437125 477396
rect 438163 477460 438229 477461
rect 438163 477396 438164 477460
rect 438228 477396 438229 477460
rect 438163 477395 438229 477396
rect 435955 477188 436021 477189
rect 435955 477124 435956 477188
rect 436020 477124 436021 477188
rect 435955 477123 436021 477124
rect 438534 477053 438594 479710
rect 439454 477189 439514 479710
rect 439451 477188 439517 477189
rect 439451 477124 439452 477188
rect 439516 477124 439517 477188
rect 439451 477123 439517 477124
rect 440742 477053 440802 479710
rect 438531 477052 438597 477053
rect 438531 476988 438532 477052
rect 438596 476988 438597 477052
rect 438531 476987 438597 476988
rect 440739 477052 440805 477053
rect 440739 476988 440740 477052
rect 440804 476988 440805 477052
rect 440739 476987 440805 476988
rect 441110 476917 441170 479710
rect 441662 479710 441820 479770
rect 442766 479710 442908 479770
rect 443502 479710 443588 479770
rect 443870 479710 443996 479770
rect 445296 479770 445356 480080
rect 445976 479770 446036 480080
rect 446384 479770 446444 480080
rect 447608 479770 447668 480080
rect 448288 479770 448348 480080
rect 448696 479770 448756 480080
rect 449784 479770 449844 480080
rect 451008 479770 451068 480080
rect 445296 479710 445402 479770
rect 441662 476917 441722 479710
rect 441107 476916 441173 476917
rect 441107 476852 441108 476916
rect 441172 476852 441173 476916
rect 441107 476851 441173 476852
rect 441659 476916 441725 476917
rect 441659 476852 441660 476916
rect 441724 476852 441725 476916
rect 441659 476851 441725 476852
rect 442766 476509 442826 479710
rect 443502 476509 443562 479710
rect 443870 477461 443930 479710
rect 443867 477460 443933 477461
rect 443867 477396 443868 477460
rect 443932 477396 443933 477460
rect 443867 477395 443933 477396
rect 445342 477189 445402 479710
rect 445894 479710 446036 479770
rect 446262 479710 446444 479770
rect 447550 479710 447668 479770
rect 448286 479710 448348 479770
rect 448654 479710 448756 479770
rect 449758 479710 449844 479770
rect 450862 479710 451068 479770
rect 445339 477188 445405 477189
rect 445339 477124 445340 477188
rect 445404 477124 445405 477188
rect 445339 477123 445405 477124
rect 433747 476508 433813 476509
rect 433747 476444 433748 476508
rect 433812 476444 433813 476508
rect 433747 476443 433813 476444
rect 442763 476508 442829 476509
rect 442763 476444 442764 476508
rect 442828 476444 442829 476508
rect 442763 476443 442829 476444
rect 443499 476508 443565 476509
rect 443499 476444 443500 476508
rect 443564 476444 443565 476508
rect 443499 476443 443565 476444
rect 445894 476237 445954 479710
rect 446262 477189 446322 479710
rect 447550 477461 447610 479710
rect 447547 477460 447613 477461
rect 447547 477396 447548 477460
rect 447612 477396 447613 477460
rect 447547 477395 447613 477396
rect 446259 477188 446325 477189
rect 446259 477124 446260 477188
rect 446324 477124 446325 477188
rect 446259 477123 446325 477124
rect 448286 476237 448346 479710
rect 448654 477189 448714 479710
rect 449758 477461 449818 479710
rect 449755 477460 449821 477461
rect 449755 477396 449756 477460
rect 449820 477396 449821 477460
rect 449755 477395 449821 477396
rect 448651 477188 448717 477189
rect 448651 477124 448652 477188
rect 448716 477124 448717 477188
rect 448651 477123 448717 477124
rect 450862 476237 450922 479710
rect 451144 479090 451204 480080
rect 452232 479770 452292 480080
rect 453320 479770 453380 480080
rect 451046 479030 451204 479090
rect 452150 479710 452292 479770
rect 453254 479710 453380 479770
rect 453592 479770 453652 480080
rect 454408 479770 454468 480080
rect 455768 479770 455828 480080
rect 456040 479770 456100 480080
rect 456992 479770 457052 480080
rect 458080 479770 458140 480080
rect 458488 479770 458548 480080
rect 459168 479770 459228 480080
rect 453592 479710 453682 479770
rect 451046 476509 451106 479030
rect 452150 477189 452210 479710
rect 453254 477461 453314 479710
rect 453251 477460 453317 477461
rect 453251 477396 453252 477460
rect 453316 477396 453317 477460
rect 453251 477395 453317 477396
rect 452147 477188 452213 477189
rect 452147 477124 452148 477188
rect 452212 477124 452213 477188
rect 452147 477123 452213 477124
rect 453622 477053 453682 479710
rect 454358 479710 454468 479770
rect 455646 479710 455828 479770
rect 456014 479710 456100 479770
rect 456934 479710 457052 479770
rect 458038 479710 458140 479770
rect 458406 479710 458548 479770
rect 459142 479710 459228 479770
rect 460936 479770 460996 480080
rect 463520 479770 463580 480080
rect 465968 479770 466028 480080
rect 468280 479770 468340 480080
rect 471000 479770 471060 480080
rect 460936 479710 461042 479770
rect 463520 479710 463618 479770
rect 454358 477053 454418 479710
rect 453619 477052 453685 477053
rect 453619 476988 453620 477052
rect 453684 476988 453685 477052
rect 453619 476987 453685 476988
rect 454355 477052 454421 477053
rect 454355 476988 454356 477052
rect 454420 476988 454421 477052
rect 454355 476987 454421 476988
rect 455646 476917 455706 479710
rect 455643 476916 455709 476917
rect 455643 476852 455644 476916
rect 455708 476852 455709 476916
rect 455643 476851 455709 476852
rect 456014 476781 456074 479710
rect 456934 477053 456994 479710
rect 456931 477052 456997 477053
rect 456931 476988 456932 477052
rect 456996 476988 456997 477052
rect 456931 476987 456997 476988
rect 458038 476917 458098 479710
rect 458035 476916 458101 476917
rect 458035 476852 458036 476916
rect 458100 476852 458101 476916
rect 458035 476851 458101 476852
rect 456011 476780 456077 476781
rect 456011 476716 456012 476780
rect 456076 476716 456077 476780
rect 456011 476715 456077 476716
rect 451043 476508 451109 476509
rect 451043 476444 451044 476508
rect 451108 476444 451109 476508
rect 451043 476443 451109 476444
rect 458406 476373 458466 479710
rect 459142 477189 459202 479710
rect 460982 477325 461042 479710
rect 460979 477324 461045 477325
rect 460979 477260 460980 477324
rect 461044 477260 461045 477324
rect 460979 477259 461045 477260
rect 463558 477189 463618 479710
rect 465950 479710 466028 479770
rect 468158 479710 468340 479770
rect 470918 479710 471060 479770
rect 473448 479770 473508 480080
rect 475896 479770 475956 480080
rect 478480 479770 478540 480080
rect 480928 479770 480988 480080
rect 483512 479770 483572 480080
rect 473448 479710 473554 479770
rect 459139 477188 459205 477189
rect 459139 477124 459140 477188
rect 459204 477124 459205 477188
rect 459139 477123 459205 477124
rect 463555 477188 463621 477189
rect 463555 477124 463556 477188
rect 463620 477124 463621 477188
rect 463555 477123 463621 477124
rect 458403 476372 458469 476373
rect 458403 476308 458404 476372
rect 458468 476308 458469 476372
rect 458403 476307 458469 476308
rect 465950 476237 466010 479710
rect 468158 476237 468218 479710
rect 470918 476237 470978 479710
rect 473494 476237 473554 479710
rect 475886 479710 475956 479770
rect 478462 479710 478540 479770
rect 480854 479710 480988 479770
rect 483430 479710 483572 479770
rect 485960 479770 486020 480080
rect 488544 479770 488604 480080
rect 490992 479770 491052 480080
rect 493440 479770 493500 480080
rect 485960 479710 486066 479770
rect 488544 479710 488642 479770
rect 475886 476509 475946 479710
rect 478462 476509 478522 479710
rect 475883 476508 475949 476509
rect 475883 476444 475884 476508
rect 475948 476444 475949 476508
rect 475883 476443 475949 476444
rect 478459 476508 478525 476509
rect 478459 476444 478460 476508
rect 478524 476444 478525 476508
rect 478459 476443 478525 476444
rect 480854 476237 480914 479710
rect 483430 476917 483490 479710
rect 483427 476916 483493 476917
rect 483427 476852 483428 476916
rect 483492 476852 483493 476916
rect 483427 476851 483493 476852
rect 486006 476237 486066 479710
rect 488582 476237 488642 479710
rect 490974 479710 491052 479770
rect 493366 479710 493500 479770
rect 495888 479770 495948 480080
rect 498472 479770 498532 480080
rect 500920 479770 500980 480080
rect 503368 479770 503428 480080
rect 505952 479770 506012 480080
rect 495888 479710 496002 479770
rect 498472 479710 498578 479770
rect 490974 476781 491034 479710
rect 490971 476780 491037 476781
rect 490971 476716 490972 476780
rect 491036 476716 491037 476780
rect 490971 476715 491037 476716
rect 493366 476237 493426 479710
rect 495942 476237 496002 479710
rect 498518 476781 498578 479710
rect 500910 479710 500980 479770
rect 503302 479710 503428 479770
rect 505878 479710 506012 479770
rect 498515 476780 498581 476781
rect 498515 476716 498516 476780
rect 498580 476716 498581 476780
rect 498515 476715 498581 476716
rect 500910 476237 500970 479710
rect 503302 476373 503362 479710
rect 503299 476372 503365 476373
rect 503299 476308 503300 476372
rect 503364 476308 503365 476372
rect 503299 476307 503365 476308
rect 505878 476237 505938 479710
rect 428227 476236 428293 476237
rect 428227 476172 428228 476236
rect 428292 476172 428293 476236
rect 428227 476171 428293 476172
rect 430619 476236 430685 476237
rect 430619 476172 430620 476236
rect 430684 476172 430685 476236
rect 430619 476171 430685 476172
rect 445891 476236 445957 476237
rect 445891 476172 445892 476236
rect 445956 476172 445957 476236
rect 445891 476171 445957 476172
rect 448283 476236 448349 476237
rect 448283 476172 448284 476236
rect 448348 476172 448349 476236
rect 448283 476171 448349 476172
rect 450859 476236 450925 476237
rect 450859 476172 450860 476236
rect 450924 476172 450925 476236
rect 450859 476171 450925 476172
rect 465947 476236 466013 476237
rect 465947 476172 465948 476236
rect 466012 476172 466013 476236
rect 465947 476171 466013 476172
rect 468155 476236 468221 476237
rect 468155 476172 468156 476236
rect 468220 476172 468221 476236
rect 468155 476171 468221 476172
rect 470915 476236 470981 476237
rect 470915 476172 470916 476236
rect 470980 476172 470981 476236
rect 470915 476171 470981 476172
rect 473491 476236 473557 476237
rect 473491 476172 473492 476236
rect 473556 476172 473557 476236
rect 473491 476171 473557 476172
rect 480851 476236 480917 476237
rect 480851 476172 480852 476236
rect 480916 476172 480917 476236
rect 480851 476171 480917 476172
rect 486003 476236 486069 476237
rect 486003 476172 486004 476236
rect 486068 476172 486069 476236
rect 486003 476171 486069 476172
rect 488579 476236 488645 476237
rect 488579 476172 488580 476236
rect 488644 476172 488645 476236
rect 488579 476171 488645 476172
rect 493363 476236 493429 476237
rect 493363 476172 493364 476236
rect 493428 476172 493429 476236
rect 493363 476171 493429 476172
rect 495939 476236 496005 476237
rect 495939 476172 495940 476236
rect 496004 476172 496005 476236
rect 495939 476171 496005 476172
rect 500907 476236 500973 476237
rect 500907 476172 500908 476236
rect 500972 476172 500973 476236
rect 500907 476171 500973 476172
rect 505875 476236 505941 476237
rect 505875 476172 505876 476236
rect 505940 476172 505941 476236
rect 505875 476171 505941 476172
rect 399523 474604 399589 474605
rect 399523 474540 399524 474604
rect 399588 474540 399589 474604
rect 399523 474539 399589 474540
rect 399526 351253 399586 474539
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 530899 446452 530965 446453
rect 530899 446388 530900 446452
rect 530964 446388 530965 446452
rect 530899 446387 530965 446388
rect 530902 443730 530962 446387
rect 530840 443670 530962 443730
rect 530840 443202 530900 443670
rect 400272 439174 400620 439206
rect 400272 438938 400328 439174
rect 400564 438938 400620 439174
rect 400272 438854 400620 438938
rect 400272 438618 400328 438854
rect 400564 438618 400620 438854
rect 400272 438586 400620 438618
rect 536000 439174 536348 439206
rect 536000 438938 536056 439174
rect 536292 438938 536348 439174
rect 536000 438854 536348 438938
rect 536000 438618 536056 438854
rect 536292 438618 536348 438854
rect 536000 438586 536348 438618
rect 400952 435454 401300 435486
rect 400952 435218 401008 435454
rect 401244 435218 401300 435454
rect 400952 435134 401300 435218
rect 400952 434898 401008 435134
rect 401244 434898 401300 435134
rect 400952 434866 401300 434898
rect 535320 435454 535668 435486
rect 535320 435218 535376 435454
rect 535612 435218 535668 435454
rect 535320 435134 535668 435218
rect 535320 434898 535376 435134
rect 535612 434898 535668 435134
rect 535320 434866 535668 434898
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 400272 403174 400620 403206
rect 400272 402938 400328 403174
rect 400564 402938 400620 403174
rect 400272 402854 400620 402938
rect 400272 402618 400328 402854
rect 400564 402618 400620 402854
rect 400272 402586 400620 402618
rect 536000 403174 536348 403206
rect 536000 402938 536056 403174
rect 536292 402938 536348 403174
rect 536000 402854 536348 402938
rect 536000 402618 536056 402854
rect 536292 402618 536348 402854
rect 536000 402586 536348 402618
rect 400952 399454 401300 399486
rect 400952 399218 401008 399454
rect 401244 399218 401300 399454
rect 400952 399134 401300 399218
rect 400952 398898 401008 399134
rect 401244 398898 401300 399134
rect 400952 398866 401300 398898
rect 535320 399454 535668 399486
rect 535320 399218 535376 399454
rect 535612 399218 535668 399454
rect 535320 399134 535668 399218
rect 535320 398898 535376 399134
rect 535612 398898 535668 399134
rect 535320 398866 535668 398898
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 400272 367174 400620 367206
rect 400272 366938 400328 367174
rect 400564 366938 400620 367174
rect 400272 366854 400620 366938
rect 400272 366618 400328 366854
rect 400564 366618 400620 366854
rect 400272 366586 400620 366618
rect 536000 367174 536348 367206
rect 536000 366938 536056 367174
rect 536292 366938 536348 367174
rect 536000 366854 536348 366938
rect 536000 366618 536056 366854
rect 536292 366618 536348 366854
rect 536000 366586 536348 366618
rect 400952 363454 401300 363486
rect 400952 363218 401008 363454
rect 401244 363218 401300 363454
rect 400952 363134 401300 363218
rect 400952 362898 401008 363134
rect 401244 362898 401300 363134
rect 400952 362866 401300 362898
rect 535320 363454 535668 363486
rect 535320 363218 535376 363454
rect 535612 363218 535668 363454
rect 535320 363134 535668 363218
rect 535320 362898 535376 363134
rect 535612 362898 535668 363134
rect 535320 362866 535668 362898
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 416056 359410 416116 360060
rect 417144 359410 417204 360060
rect 418232 359410 418292 360060
rect 419592 359410 419652 360060
rect 420544 359410 420604 360060
rect 416056 359350 416146 359410
rect 417144 359350 417250 359410
rect 416086 358189 416146 359350
rect 416083 358188 416149 358189
rect 416083 358124 416084 358188
rect 416148 358124 416149 358188
rect 416083 358123 416149 358124
rect 399523 351252 399589 351253
rect 399523 351188 399524 351252
rect 399588 351188 399589 351252
rect 399523 351187 399589 351188
rect 399339 348396 399405 348397
rect 399339 348332 399340 348396
rect 399404 348332 399405 348396
rect 399339 348331 399405 348332
rect 401514 331174 402134 358064
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 398787 311132 398853 311133
rect 398787 311068 398788 311132
rect 398852 311068 398853 311132
rect 398787 311067 398853 311068
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 394928 219454 395248 219486
rect 394928 219218 394970 219454
rect 395206 219218 395248 219454
rect 394928 219134 395248 219218
rect 394928 218898 394970 219134
rect 395206 218898 395248 219134
rect 394928 218866 395248 218898
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 394928 183454 395248 183486
rect 394928 183218 394970 183454
rect 395206 183218 395248 183454
rect 394928 183134 395248 183218
rect 394928 182898 394970 183134
rect 395206 182898 395248 183134
rect 394928 182866 395248 182898
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 394928 147454 395248 147486
rect 394928 147218 394970 147454
rect 395206 147218 395248 147454
rect 394928 147134 395248 147218
rect 394928 146898 394970 147134
rect 395206 146898 395248 147134
rect 394928 146866 395248 146898
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 394928 111454 395248 111486
rect 394928 111218 394970 111454
rect 395206 111218 395248 111454
rect 394928 111134 395248 111218
rect 394928 110898 394970 111134
rect 395206 110898 395248 111134
rect 394928 110866 395248 110898
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 394928 75454 395248 75486
rect 394928 75218 394970 75454
rect 395206 75218 395248 75454
rect 394928 75134 395248 75218
rect 394928 74898 394970 75134
rect 395206 74898 395248 75134
rect 394928 74866 395248 74898
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 405234 334894 405854 358064
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 228961 405854 262338
rect 408954 338614 409574 358064
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 228961 409574 230058
rect 412674 342334 413294 358064
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 306334 413294 341778
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 228961 413294 233778
rect 416394 346054 417014 358064
rect 417190 357373 417250 359350
rect 418110 359350 418292 359410
rect 419582 359350 419652 359410
rect 419950 359350 420604 359410
rect 421768 359410 421828 360060
rect 423128 359410 423188 360060
rect 421768 359350 421850 359410
rect 417187 357372 417253 357373
rect 417187 357308 417188 357372
rect 417252 357308 417253 357372
rect 417187 357307 417253 357308
rect 418110 357237 418170 359350
rect 418107 357236 418173 357237
rect 418107 357172 418108 357236
rect 418172 357172 418173 357236
rect 418107 357171 418173 357172
rect 419582 357101 419642 359350
rect 419579 357100 419645 357101
rect 419579 357036 419580 357100
rect 419644 357036 419645 357100
rect 419579 357035 419645 357036
rect 419950 356965 420010 359350
rect 419947 356964 420013 356965
rect 419947 356900 419948 356964
rect 420012 356900 420013 356964
rect 419947 356899 420013 356900
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 416394 310054 417014 345498
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 228961 417014 237498
rect 420114 349774 420734 357940
rect 421790 356829 421850 359350
rect 423078 359350 423188 359410
rect 424216 359410 424276 360060
rect 425440 359410 425500 360060
rect 426528 359410 426588 360060
rect 427616 359410 427676 360060
rect 428296 359410 428356 360060
rect 428704 359410 428764 360060
rect 424216 359350 424610 359410
rect 425440 359350 425530 359410
rect 426528 359350 426634 359410
rect 427616 359350 427738 359410
rect 423078 357373 423138 359350
rect 423075 357372 423141 357373
rect 423075 357308 423076 357372
rect 423140 357308 423141 357372
rect 423075 357307 423141 357308
rect 421787 356828 421853 356829
rect 421787 356764 421788 356828
rect 421852 356764 421853 356828
rect 421787 356763 421853 356764
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 420114 313774 420734 349218
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 228961 420734 241218
rect 423834 353494 424454 357940
rect 424550 357373 424610 359350
rect 425470 357373 425530 359350
rect 426574 357373 426634 359350
rect 427678 357373 427738 359350
rect 428230 359350 428356 359410
rect 428598 359350 428764 359410
rect 430064 359410 430124 360060
rect 430744 359410 430804 360060
rect 431288 359410 431348 360060
rect 432376 359410 432436 360060
rect 433464 359410 433524 360060
rect 430064 359350 430130 359410
rect 428230 357373 428290 359350
rect 428598 357373 428658 359350
rect 430070 357373 430130 359350
rect 430622 359350 430804 359410
rect 431174 359350 431348 359410
rect 431726 359350 432436 359410
rect 433382 359350 433524 359410
rect 433600 359410 433660 360060
rect 434552 359410 434612 360060
rect 435912 359410 435972 360060
rect 433600 359350 433810 359410
rect 434552 359350 434730 359410
rect 430622 357373 430682 359350
rect 424547 357372 424613 357373
rect 424547 357308 424548 357372
rect 424612 357308 424613 357372
rect 424547 357307 424613 357308
rect 425467 357372 425533 357373
rect 425467 357308 425468 357372
rect 425532 357308 425533 357372
rect 425467 357307 425533 357308
rect 426571 357372 426637 357373
rect 426571 357308 426572 357372
rect 426636 357308 426637 357372
rect 426571 357307 426637 357308
rect 427675 357372 427741 357373
rect 427675 357308 427676 357372
rect 427740 357308 427741 357372
rect 427675 357307 427741 357308
rect 428227 357372 428293 357373
rect 428227 357308 428228 357372
rect 428292 357308 428293 357372
rect 428227 357307 428293 357308
rect 428595 357372 428661 357373
rect 428595 357308 428596 357372
rect 428660 357308 428661 357372
rect 428595 357307 428661 357308
rect 430067 357372 430133 357373
rect 430067 357308 430068 357372
rect 430132 357308 430133 357372
rect 430067 357307 430133 357308
rect 430619 357372 430685 357373
rect 430619 357308 430620 357372
rect 430684 357308 430685 357372
rect 430619 357307 430685 357308
rect 431174 357237 431234 359350
rect 431726 357370 431786 359350
rect 431907 357372 431973 357373
rect 431907 357370 431908 357372
rect 431726 357310 431908 357370
rect 431907 357308 431908 357310
rect 431972 357308 431973 357372
rect 431907 357307 431973 357308
rect 433382 357237 433442 359350
rect 433750 358730 433810 359350
rect 433566 358670 433810 358730
rect 433566 357373 433626 358670
rect 433563 357372 433629 357373
rect 433563 357308 433564 357372
rect 433628 357308 433629 357372
rect 433563 357307 433629 357308
rect 431171 357236 431237 357237
rect 431171 357172 431172 357236
rect 431236 357172 431237 357236
rect 431171 357171 431237 357172
rect 433379 357236 433445 357237
rect 433379 357172 433380 357236
rect 433444 357172 433445 357236
rect 433379 357171 433445 357172
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 423834 317494 424454 352938
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 228961 424454 244938
rect 433794 327454 434414 358064
rect 434670 357237 434730 359350
rect 435774 359350 435972 359410
rect 435774 357237 435834 359350
rect 436048 358730 436108 360060
rect 437000 359410 437060 360060
rect 438088 359410 438148 360060
rect 438496 359410 438556 360060
rect 439448 359410 439508 360060
rect 440672 359410 440732 360060
rect 441080 359410 441140 360060
rect 437000 359350 437122 359410
rect 438088 359350 438410 359410
rect 438496 359350 438594 359410
rect 439448 359350 439514 359410
rect 440672 359350 440802 359410
rect 435958 358670 436108 358730
rect 435958 357373 436018 358670
rect 437062 357373 437122 359350
rect 435955 357372 436021 357373
rect 435955 357308 435956 357372
rect 436020 357308 436021 357372
rect 435955 357307 436021 357308
rect 437059 357372 437125 357373
rect 437059 357308 437060 357372
rect 437124 357308 437125 357372
rect 437059 357307 437125 357308
rect 434667 357236 434733 357237
rect 434667 357172 434668 357236
rect 434732 357172 434733 357236
rect 434667 357171 434733 357172
rect 435771 357236 435837 357237
rect 435771 357172 435772 357236
rect 435836 357172 435837 357236
rect 435771 357171 435837 357172
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 228961 434414 254898
rect 437514 331174 438134 357940
rect 438350 357237 438410 359350
rect 438534 357373 438594 359350
rect 438531 357372 438597 357373
rect 438531 357308 438532 357372
rect 438596 357308 438597 357372
rect 438531 357307 438597 357308
rect 439454 357237 439514 359350
rect 438347 357236 438413 357237
rect 438347 357172 438348 357236
rect 438412 357172 438413 357236
rect 438347 357171 438413 357172
rect 438899 357236 438965 357237
rect 438899 357172 438900 357236
rect 438964 357172 438965 357236
rect 438899 357171 438965 357172
rect 439451 357236 439517 357237
rect 439451 357172 439452 357236
rect 439516 357172 439517 357236
rect 439451 357171 439517 357172
rect 438902 356421 438962 357171
rect 440742 356557 440802 359350
rect 440926 359350 441140 359410
rect 441760 359410 441820 360060
rect 442848 359410 442908 360060
rect 443528 359410 443588 360060
rect 443936 359410 443996 360060
rect 445296 359410 445356 360060
rect 445976 359410 446036 360060
rect 446384 359410 446444 360060
rect 447608 359410 447668 360060
rect 448288 359410 448348 360060
rect 448696 359410 448756 360060
rect 449784 359410 449844 360060
rect 450859 359548 450925 359549
rect 450859 359484 450860 359548
rect 450924 359484 450925 359548
rect 450859 359483 450925 359484
rect 441760 359350 442090 359410
rect 440926 357373 440986 359350
rect 440923 357372 440989 357373
rect 440923 357308 440924 357372
rect 440988 357308 440989 357372
rect 440923 357307 440989 357308
rect 440739 356556 440805 356557
rect 440739 356492 440740 356556
rect 440804 356492 440805 356556
rect 440739 356491 440805 356492
rect 438899 356420 438965 356421
rect 438899 356356 438900 356420
rect 438964 356356 438965 356420
rect 438899 356355 438965 356356
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 228961 438134 258618
rect 441234 334894 441854 357940
rect 442030 356557 442090 359350
rect 442766 359350 442908 359410
rect 443502 359350 443588 359410
rect 443870 359350 443996 359410
rect 444790 359350 445356 359410
rect 445894 359350 446036 359410
rect 446262 359350 446444 359410
rect 447550 359350 447668 359410
rect 448286 359350 448348 359410
rect 448470 359350 448756 359410
rect 449758 359350 449844 359410
rect 442027 356556 442093 356557
rect 442027 356492 442028 356556
rect 442092 356492 442093 356556
rect 442027 356491 442093 356492
rect 442766 356421 442826 359350
rect 443502 357237 443562 359350
rect 443499 357236 443565 357237
rect 443499 357172 443500 357236
rect 443564 357172 443565 357236
rect 443499 357171 443565 357172
rect 443870 356557 443930 359350
rect 443867 356556 443933 356557
rect 443867 356492 443868 356556
rect 443932 356492 443933 356556
rect 443867 356491 443933 356492
rect 444790 356421 444850 359350
rect 442763 356420 442829 356421
rect 442763 356356 442764 356420
rect 442828 356356 442829 356420
rect 442763 356355 442829 356356
rect 444787 356420 444853 356421
rect 444787 356356 444788 356420
rect 444852 356356 444853 356420
rect 444787 356355 444853 356356
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 229452 441854 262338
rect 444954 338614 445574 357940
rect 445894 357373 445954 359350
rect 445891 357372 445957 357373
rect 445891 357308 445892 357372
rect 445956 357308 445957 357372
rect 445891 357307 445957 357308
rect 446262 356693 446322 359350
rect 447550 357101 447610 359350
rect 448286 357373 448346 359350
rect 448283 357372 448349 357373
rect 448283 357308 448284 357372
rect 448348 357308 448349 357372
rect 448283 357307 448349 357308
rect 447547 357100 447613 357101
rect 447547 357036 447548 357100
rect 447612 357036 447613 357100
rect 447547 357035 447613 357036
rect 448470 356829 448530 359350
rect 448467 356828 448533 356829
rect 448467 356764 448468 356828
rect 448532 356764 448533 356828
rect 448467 356763 448533 356764
rect 446259 356692 446325 356693
rect 446259 356628 446260 356692
rect 446324 356628 446325 356692
rect 446259 356627 446325 356628
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 228961 445574 230058
rect 448674 342334 449294 357940
rect 449758 356557 449818 359350
rect 450862 357101 450922 359483
rect 451008 359410 451068 360060
rect 451144 359549 451204 360060
rect 451141 359548 451207 359549
rect 451141 359484 451142 359548
rect 451206 359484 451207 359548
rect 452232 359546 452292 360060
rect 453320 359546 453380 360060
rect 451141 359483 451207 359484
rect 452150 359486 452292 359546
rect 453254 359486 453380 359546
rect 453592 359546 453652 360060
rect 454408 359546 454468 360060
rect 455768 359546 455828 360060
rect 456040 359546 456100 360060
rect 456992 359546 457052 360060
rect 458080 359546 458140 360060
rect 458488 359546 458548 360060
rect 459168 359546 459228 360060
rect 453592 359486 453682 359546
rect 451008 359350 451106 359410
rect 451046 357373 451106 359350
rect 452150 357373 452210 359486
rect 451043 357372 451109 357373
rect 451043 357308 451044 357372
rect 451108 357308 451109 357372
rect 451043 357307 451109 357308
rect 452147 357372 452213 357373
rect 452147 357308 452148 357372
rect 452212 357308 452213 357372
rect 452147 357307 452213 357308
rect 450859 357100 450925 357101
rect 450859 357036 450860 357100
rect 450924 357036 450925 357100
rect 450859 357035 450925 357036
rect 449755 356556 449821 356557
rect 449755 356492 449756 356556
rect 449820 356492 449821 356556
rect 449755 356491 449821 356492
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448674 306334 449294 341778
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 228961 449294 233778
rect 452394 346054 453014 358064
rect 453254 356965 453314 359486
rect 453622 357373 453682 359486
rect 454358 359486 454468 359546
rect 455646 359486 455828 359546
rect 456014 359486 456100 359546
rect 456934 359486 457052 359546
rect 458038 359486 458140 359546
rect 458406 359486 458548 359546
rect 459142 359486 459228 359546
rect 453619 357372 453685 357373
rect 453619 357308 453620 357372
rect 453684 357308 453685 357372
rect 453619 357307 453685 357308
rect 454358 357101 454418 359486
rect 454355 357100 454421 357101
rect 454355 357036 454356 357100
rect 454420 357036 454421 357100
rect 454355 357035 454421 357036
rect 455646 356965 455706 359486
rect 456014 358730 456074 359486
rect 455830 358670 456074 358730
rect 455830 357373 455890 358670
rect 455827 357372 455893 357373
rect 455827 357308 455828 357372
rect 455892 357308 455893 357372
rect 455827 357307 455893 357308
rect 453251 356964 453317 356965
rect 453251 356900 453252 356964
rect 453316 356900 453317 356964
rect 453251 356899 453317 356900
rect 455643 356964 455709 356965
rect 455643 356900 455644 356964
rect 455708 356900 455709 356964
rect 455643 356899 455709 356900
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 452394 310054 453014 345498
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 228961 453014 237498
rect 456114 349774 456734 357940
rect 456934 356829 456994 359486
rect 458038 357237 458098 359486
rect 458406 357373 458466 359486
rect 458403 357372 458469 357373
rect 458403 357308 458404 357372
rect 458468 357308 458469 357372
rect 458403 357307 458469 357308
rect 459142 357237 459202 359486
rect 460936 359410 460996 360060
rect 463520 359410 463580 360060
rect 465968 359410 466028 360060
rect 468280 359410 468340 360060
rect 471000 359410 471060 360060
rect 473448 359410 473508 360060
rect 475896 359410 475956 360060
rect 478480 359410 478540 360060
rect 480928 359410 480988 360060
rect 483512 359410 483572 360060
rect 460936 359350 461042 359410
rect 463520 359350 463618 359410
rect 458035 357236 458101 357237
rect 458035 357172 458036 357236
rect 458100 357172 458101 357236
rect 458035 357171 458101 357172
rect 459139 357236 459205 357237
rect 459139 357172 459140 357236
rect 459204 357172 459205 357236
rect 459139 357171 459205 357172
rect 456931 356828 456997 356829
rect 456931 356764 456932 356828
rect 456996 356764 456997 356828
rect 456931 356763 456997 356764
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 229452 456734 241218
rect 459834 353494 460454 358064
rect 460982 356149 461042 359350
rect 463558 357373 463618 359350
rect 465950 359350 466028 359410
rect 468158 359350 468340 359410
rect 470918 359350 471060 359410
rect 473310 359350 473508 359410
rect 475886 359350 475956 359410
rect 478462 359350 478540 359410
rect 480670 359350 480988 359410
rect 483430 359350 483572 359410
rect 485960 359410 486020 360060
rect 488544 359410 488604 360060
rect 490992 359410 491052 360060
rect 493440 359410 493500 360060
rect 495888 359410 495948 360060
rect 485960 359350 486066 359410
rect 488544 359350 488642 359410
rect 465950 357373 466010 359350
rect 468158 357373 468218 359350
rect 463555 357372 463621 357373
rect 463555 357308 463556 357372
rect 463620 357308 463621 357372
rect 463555 357307 463621 357308
rect 465947 357372 466013 357373
rect 465947 357308 465948 357372
rect 466012 357308 466013 357372
rect 465947 357307 466013 357308
rect 468155 357372 468221 357373
rect 468155 357308 468156 357372
rect 468220 357308 468221 357372
rect 468155 357307 468221 357308
rect 460979 356148 461045 356149
rect 460979 356084 460980 356148
rect 461044 356084 461045 356148
rect 460979 356083 461045 356084
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 228961 460454 244938
rect 469794 327454 470414 358064
rect 470918 356285 470978 359350
rect 473310 357373 473370 359350
rect 473307 357372 473373 357373
rect 473307 357308 473308 357372
rect 473372 357308 473373 357372
rect 473307 357307 473373 357308
rect 470915 356284 470981 356285
rect 470915 356220 470916 356284
rect 470980 356220 470981 356284
rect 470915 356219 470981 356220
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 228961 470414 254898
rect 473514 331174 474134 357940
rect 475886 356421 475946 359350
rect 475883 356420 475949 356421
rect 475883 356356 475884 356420
rect 475948 356356 475949 356420
rect 475883 356355 475949 356356
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 228961 474134 258618
rect 477234 334894 477854 358064
rect 478462 357373 478522 359350
rect 478459 357372 478525 357373
rect 478459 357308 478460 357372
rect 478524 357308 478525 357372
rect 478459 357307 478525 357308
rect 480670 357101 480730 359350
rect 480667 357100 480733 357101
rect 480667 357036 480668 357100
rect 480732 357036 480733 357100
rect 480667 357035 480733 357036
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 228961 477854 262338
rect 480954 338614 481574 357940
rect 483430 356557 483490 359350
rect 483427 356556 483493 356557
rect 483427 356492 483428 356556
rect 483492 356492 483493 356556
rect 483427 356491 483493 356492
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 228961 481574 230058
rect 484674 342334 485294 358064
rect 486006 357373 486066 359350
rect 488582 358189 488642 359350
rect 489686 359350 491052 359410
rect 493366 359350 493500 359410
rect 495574 359350 495948 359410
rect 498472 359410 498532 360060
rect 500920 359410 500980 360060
rect 503368 359410 503428 360060
rect 505952 359410 506012 360060
rect 498472 359350 498578 359410
rect 488579 358188 488645 358189
rect 488579 358124 488580 358188
rect 488644 358124 488645 358188
rect 488579 358123 488645 358124
rect 486003 357372 486069 357373
rect 486003 357308 486004 357372
rect 486068 357308 486069 357372
rect 486003 357307 486069 357308
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 484674 306334 485294 341778
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 234334 485294 269778
rect 484674 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 485294 234334
rect 484674 234014 485294 234098
rect 484674 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 485294 234014
rect 484674 228961 485294 233778
rect 488394 346054 489014 357940
rect 489686 356285 489746 359350
rect 489683 356284 489749 356285
rect 489683 356220 489684 356284
rect 489748 356220 489749 356284
rect 489683 356219 489749 356220
rect 488394 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 489014 346054
rect 488394 345734 489014 345818
rect 488394 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 489014 345734
rect 488394 310054 489014 345498
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 238054 489014 273498
rect 488394 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 489014 238054
rect 488394 237734 489014 237818
rect 488394 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 489014 237734
rect 488394 228961 489014 237498
rect 492114 349774 492734 358064
rect 493366 356149 493426 359350
rect 495574 356285 495634 359350
rect 495571 356284 495637 356285
rect 495571 356220 495572 356284
rect 495636 356220 495637 356284
rect 495571 356219 495637 356220
rect 493363 356148 493429 356149
rect 493363 356084 493364 356148
rect 493428 356084 493429 356148
rect 493363 356083 493429 356084
rect 492114 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 492734 349774
rect 492114 349454 492734 349538
rect 492114 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 492734 349454
rect 492114 313774 492734 349218
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 241774 492734 277218
rect 492114 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 492734 241774
rect 492114 241454 492734 241538
rect 492114 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 492734 241454
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 410288 223174 410608 223206
rect 410288 222938 410330 223174
rect 410566 222938 410608 223174
rect 410288 222854 410608 222938
rect 410288 222618 410330 222854
rect 410566 222618 410608 222854
rect 410288 222586 410608 222618
rect 441008 223174 441328 223206
rect 441008 222938 441050 223174
rect 441286 222938 441328 223174
rect 441008 222854 441328 222938
rect 441008 222618 441050 222854
rect 441286 222618 441328 222854
rect 441008 222586 441328 222618
rect 471728 223174 472048 223206
rect 471728 222938 471770 223174
rect 472006 222938 472048 223174
rect 471728 222854 472048 222938
rect 471728 222618 471770 222854
rect 472006 222618 472048 222854
rect 471728 222586 472048 222618
rect 425648 219454 425968 219486
rect 425648 219218 425690 219454
rect 425926 219218 425968 219454
rect 425648 219134 425968 219218
rect 425648 218898 425690 219134
rect 425926 218898 425968 219134
rect 425648 218866 425968 218898
rect 456368 219454 456688 219486
rect 456368 219218 456410 219454
rect 456646 219218 456688 219454
rect 456368 219134 456688 219218
rect 456368 218898 456410 219134
rect 456646 218898 456688 219134
rect 456368 218866 456688 218898
rect 487088 219454 487408 219486
rect 487088 219218 487130 219454
rect 487366 219218 487408 219454
rect 487088 219134 487408 219218
rect 487088 218898 487130 219134
rect 487366 218898 487408 219134
rect 487088 218866 487408 218898
rect 492114 205774 492734 241218
rect 492114 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 492734 205774
rect 492114 205454 492734 205538
rect 492114 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 492734 205454
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 410288 187174 410608 187206
rect 410288 186938 410330 187174
rect 410566 186938 410608 187174
rect 410288 186854 410608 186938
rect 410288 186618 410330 186854
rect 410566 186618 410608 186854
rect 410288 186586 410608 186618
rect 441008 187174 441328 187206
rect 441008 186938 441050 187174
rect 441286 186938 441328 187174
rect 441008 186854 441328 186938
rect 441008 186618 441050 186854
rect 441286 186618 441328 186854
rect 441008 186586 441328 186618
rect 471728 187174 472048 187206
rect 471728 186938 471770 187174
rect 472006 186938 472048 187174
rect 471728 186854 472048 186938
rect 471728 186618 471770 186854
rect 472006 186618 472048 186854
rect 471728 186586 472048 186618
rect 425648 183454 425968 183486
rect 425648 183218 425690 183454
rect 425926 183218 425968 183454
rect 425648 183134 425968 183218
rect 425648 182898 425690 183134
rect 425926 182898 425968 183134
rect 425648 182866 425968 182898
rect 456368 183454 456688 183486
rect 456368 183218 456410 183454
rect 456646 183218 456688 183454
rect 456368 183134 456688 183218
rect 456368 182898 456410 183134
rect 456646 182898 456688 183134
rect 456368 182866 456688 182898
rect 487088 183454 487408 183486
rect 487088 183218 487130 183454
rect 487366 183218 487408 183454
rect 487088 183134 487408 183218
rect 487088 182898 487130 183134
rect 487366 182898 487408 183134
rect 487088 182866 487408 182898
rect 492114 169774 492734 205218
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 410288 151174 410608 151206
rect 410288 150938 410330 151174
rect 410566 150938 410608 151174
rect 410288 150854 410608 150938
rect 410288 150618 410330 150854
rect 410566 150618 410608 150854
rect 410288 150586 410608 150618
rect 441008 151174 441328 151206
rect 441008 150938 441050 151174
rect 441286 150938 441328 151174
rect 441008 150854 441328 150938
rect 441008 150618 441050 150854
rect 441286 150618 441328 150854
rect 441008 150586 441328 150618
rect 471728 151174 472048 151206
rect 471728 150938 471770 151174
rect 472006 150938 472048 151174
rect 471728 150854 472048 150938
rect 471728 150618 471770 150854
rect 472006 150618 472048 150854
rect 471728 150586 472048 150618
rect 425648 147454 425968 147486
rect 425648 147218 425690 147454
rect 425926 147218 425968 147454
rect 425648 147134 425968 147218
rect 425648 146898 425690 147134
rect 425926 146898 425968 147134
rect 425648 146866 425968 146898
rect 456368 147454 456688 147486
rect 456368 147218 456410 147454
rect 456646 147218 456688 147454
rect 456368 147134 456688 147218
rect 456368 146898 456410 147134
rect 456646 146898 456688 147134
rect 456368 146866 456688 146898
rect 487088 147454 487408 147486
rect 487088 147218 487130 147454
rect 487366 147218 487408 147454
rect 487088 147134 487408 147218
rect 487088 146898 487130 147134
rect 487366 146898 487408 147134
rect 487088 146866 487408 146898
rect 492114 133774 492734 169218
rect 492114 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 492734 133774
rect 492114 133454 492734 133538
rect 492114 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 492734 133454
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 410288 115174 410608 115206
rect 410288 114938 410330 115174
rect 410566 114938 410608 115174
rect 410288 114854 410608 114938
rect 410288 114618 410330 114854
rect 410566 114618 410608 114854
rect 410288 114586 410608 114618
rect 441008 115174 441328 115206
rect 441008 114938 441050 115174
rect 441286 114938 441328 115174
rect 441008 114854 441328 114938
rect 441008 114618 441050 114854
rect 441286 114618 441328 114854
rect 441008 114586 441328 114618
rect 471728 115174 472048 115206
rect 471728 114938 471770 115174
rect 472006 114938 472048 115174
rect 471728 114854 472048 114938
rect 471728 114618 471770 114854
rect 472006 114618 472048 114854
rect 471728 114586 472048 114618
rect 425648 111454 425968 111486
rect 425648 111218 425690 111454
rect 425926 111218 425968 111454
rect 425648 111134 425968 111218
rect 425648 110898 425690 111134
rect 425926 110898 425968 111134
rect 425648 110866 425968 110898
rect 456368 111454 456688 111486
rect 456368 111218 456410 111454
rect 456646 111218 456688 111454
rect 456368 111134 456688 111218
rect 456368 110898 456410 111134
rect 456646 110898 456688 111134
rect 456368 110866 456688 110898
rect 487088 111454 487408 111486
rect 487088 111218 487130 111454
rect 487366 111218 487408 111454
rect 487088 111134 487408 111218
rect 487088 110898 487130 111134
rect 487366 110898 487408 111134
rect 487088 110866 487408 110898
rect 492114 97774 492734 133218
rect 492114 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 492734 97774
rect 492114 97454 492734 97538
rect 492114 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 492734 97454
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 410288 79174 410608 79206
rect 410288 78938 410330 79174
rect 410566 78938 410608 79174
rect 410288 78854 410608 78938
rect 410288 78618 410330 78854
rect 410566 78618 410608 78854
rect 410288 78586 410608 78618
rect 441008 79174 441328 79206
rect 441008 78938 441050 79174
rect 441286 78938 441328 79174
rect 441008 78854 441328 78938
rect 441008 78618 441050 78854
rect 441286 78618 441328 78854
rect 441008 78586 441328 78618
rect 471728 79174 472048 79206
rect 471728 78938 471770 79174
rect 472006 78938 472048 79174
rect 471728 78854 472048 78938
rect 471728 78618 471770 78854
rect 472006 78618 472048 78854
rect 471728 78586 472048 78618
rect 425648 75454 425968 75486
rect 425648 75218 425690 75454
rect 425926 75218 425968 75454
rect 425648 75134 425968 75218
rect 425648 74898 425690 75134
rect 425926 74898 425968 75134
rect 425648 74866 425968 74898
rect 456368 75454 456688 75486
rect 456368 75218 456410 75454
rect 456646 75218 456688 75454
rect 456368 75134 456688 75218
rect 456368 74898 456410 75134
rect 456646 74898 456688 75134
rect 456368 74866 456688 74898
rect 487088 75454 487408 75486
rect 487088 75218 487130 75454
rect 487366 75218 487408 75454
rect 487088 75134 487408 75218
rect 487088 74898 487130 75134
rect 487366 74898 487408 75134
rect 487088 74866 487408 74898
rect 492114 61774 492734 97218
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 46894 405854 51375
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 50614 409574 51375
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 18334 413294 51375
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 51375
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 25774 420734 51375
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 29494 424454 51375
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 39454 434414 51375
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 43174 438134 51375
rect 444954 50614 445574 51375
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 46894 441854 50068
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 51375
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 51375
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 25774 456734 50068
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 51375
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 39454 470414 51375
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 43174 474134 51375
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 46894 477854 51375
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 50614 481574 51375
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 18334 485294 51375
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 22054 489014 51375
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 353494 496454 357940
rect 498518 357373 498578 359350
rect 500910 359350 500980 359410
rect 503302 359350 503428 359410
rect 505510 359350 506012 359410
rect 498515 357372 498581 357373
rect 498515 357308 498516 357372
rect 498580 357308 498581 357372
rect 498515 357307 498581 357308
rect 500910 356421 500970 359350
rect 503302 356829 503362 359350
rect 503299 356828 503365 356829
rect 503299 356764 503300 356828
rect 503364 356764 503365 356828
rect 503299 356763 503365 356764
rect 500907 356420 500973 356421
rect 500907 356356 500908 356420
rect 500972 356356 500973 356420
rect 500907 356355 500973 356356
rect 505510 356149 505570 359350
rect 505507 356148 505573 356149
rect 505507 356084 505508 356148
rect 505572 356084 505573 356148
rect 505507 356083 505573 356084
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 495834 317494 496454 352938
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 245494 496454 280938
rect 495834 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 496454 245494
rect 495834 245174 496454 245258
rect 495834 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 496454 245174
rect 495834 209494 496454 244938
rect 505794 327454 506414 357940
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 502448 223174 502768 223206
rect 502448 222938 502490 223174
rect 502726 222938 502768 223174
rect 502448 222854 502768 222938
rect 502448 222618 502490 222854
rect 502726 222618 502768 222854
rect 502448 222586 502768 222618
rect 495834 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 496454 209494
rect 495834 209174 496454 209258
rect 495834 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 496454 209174
rect 495834 173494 496454 208938
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 502448 187174 502768 187206
rect 502448 186938 502490 187174
rect 502726 186938 502768 187174
rect 502448 186854 502768 186938
rect 502448 186618 502490 186854
rect 502726 186618 502768 186854
rect 502448 186586 502768 186618
rect 495834 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 496454 173494
rect 495834 173174 496454 173258
rect 495834 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 496454 173174
rect 495834 137494 496454 172938
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 502448 151174 502768 151206
rect 502448 150938 502490 151174
rect 502726 150938 502768 151174
rect 502448 150854 502768 150938
rect 502448 150618 502490 150854
rect 502726 150618 502768 150854
rect 502448 150586 502768 150618
rect 495834 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 496454 137494
rect 495834 137174 496454 137258
rect 495834 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 496454 137174
rect 495834 101494 496454 136938
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 502448 115174 502768 115206
rect 502448 114938 502490 115174
rect 502726 114938 502768 115174
rect 502448 114854 502768 114938
rect 502448 114618 502490 114854
rect 502726 114618 502768 114854
rect 502448 114586 502768 114618
rect 495834 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 496454 101494
rect 495834 101174 496454 101258
rect 495834 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 496454 101174
rect 495834 65494 496454 100938
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 502448 79174 502768 79206
rect 502448 78938 502490 79174
rect 502726 78938 502768 79174
rect 502448 78854 502768 78938
rect 502448 78618 502490 78854
rect 502726 78618 502768 78854
rect 502448 78586 502768 78618
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 331174 510134 358064
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 334894 513854 358064
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 338614 517574 358064
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 520674 342334 521294 358064
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 517808 219454 518128 219486
rect 517808 219218 517850 219454
rect 518086 219218 518128 219454
rect 517808 219134 518128 219218
rect 517808 218898 517850 219134
rect 518086 218898 518128 219134
rect 517808 218866 518128 218898
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 517808 183454 518128 183486
rect 517808 183218 517850 183454
rect 518086 183218 518128 183454
rect 517808 183134 518128 183218
rect 517808 182898 517850 183134
rect 518086 182898 518128 183134
rect 517808 182866 518128 182898
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 517808 147454 518128 147486
rect 517808 147218 517850 147454
rect 518086 147218 518128 147454
rect 517808 147134 518128 147218
rect 517808 146898 517850 147134
rect 518086 146898 518128 147134
rect 517808 146866 518128 146898
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 520674 126334 521294 161778
rect 520674 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 521294 126334
rect 520674 126014 521294 126098
rect 520674 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 521294 126014
rect 517808 111454 518128 111486
rect 517808 111218 517850 111454
rect 518086 111218 518128 111454
rect 517808 111134 518128 111218
rect 517808 110898 517850 111134
rect 518086 110898 518128 111134
rect 517808 110866 518128 110898
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 520674 90334 521294 125778
rect 520674 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 521294 90334
rect 520674 90014 521294 90098
rect 520674 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 521294 90014
rect 517808 75454 518128 75486
rect 517808 75218 517850 75454
rect 518086 75218 518128 75454
rect 517808 75134 518128 75218
rect 517808 74898 517850 75134
rect 518086 74898 518128 75134
rect 517808 74866 518128 74898
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 89778
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 346054 525014 358064
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 166054 525014 201498
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 130054 525014 165498
rect 524394 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 525014 130054
rect 524394 129734 525014 129818
rect 524394 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 525014 129734
rect 524394 94054 525014 129498
rect 524394 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 525014 94054
rect 524394 93734 525014 93818
rect 524394 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 525014 93734
rect 524394 58054 525014 93498
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 349774 528734 358064
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 169774 528734 205218
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 133774 528734 169218
rect 528114 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 528734 133774
rect 528114 133454 528734 133538
rect 528114 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 528734 133454
rect 528114 97774 528734 133218
rect 528114 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 528734 97774
rect 528114 97454 528734 97538
rect 528114 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 528734 97454
rect 528114 61774 528734 97218
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 353494 532454 358064
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 533168 223174 533488 223206
rect 533168 222938 533210 223174
rect 533446 222938 533488 223174
rect 533168 222854 533488 222938
rect 533168 222618 533210 222854
rect 533446 222618 533488 222854
rect 533168 222586 533488 222618
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 173494 532454 208938
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 533168 187174 533488 187206
rect 533168 186938 533210 187174
rect 533446 186938 533488 187174
rect 533168 186854 533488 186938
rect 533168 186618 533210 186854
rect 533446 186618 533488 186854
rect 533168 186586 533488 186618
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 533168 151174 533488 151206
rect 533168 150938 533210 151174
rect 533446 150938 533488 151174
rect 533168 150854 533488 150938
rect 533168 150618 533210 150854
rect 533446 150618 533488 150854
rect 533168 150586 533488 150618
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 533168 115174 533488 115206
rect 533168 114938 533210 115174
rect 533446 114938 533488 115174
rect 533168 114854 533488 114938
rect 533168 114618 533210 114854
rect 533446 114618 533488 114854
rect 533168 114586 533488 114618
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 533168 79174 533488 79206
rect 533168 78938 533210 79174
rect 533446 78938 533488 79174
rect 533168 78854 533488 78938
rect 533168 78618 533210 78854
rect 533446 78618 533488 78854
rect 533168 78586 533488 78618
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 40328 654938 40564 655174
rect 40328 654618 40564 654854
rect 176056 654938 176292 655174
rect 176056 654618 176292 654854
rect 41008 651218 41244 651454
rect 41008 650898 41244 651134
rect 175376 651218 175612 651454
rect 175376 650898 175612 651134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 40328 618938 40564 619174
rect 40328 618618 40564 618854
rect 176056 618938 176292 619174
rect 176056 618618 176292 618854
rect 41008 615218 41244 615454
rect 41008 614898 41244 615134
rect 175376 615218 175612 615454
rect 175376 614898 175612 615134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 40328 546938 40564 547174
rect 40328 546618 40564 546854
rect 176056 546938 176292 547174
rect 176056 546618 176292 546854
rect 41008 543218 41244 543454
rect 41008 542898 41244 543134
rect 175376 543218 175612 543454
rect 175376 542898 175612 543134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 40328 510938 40564 511174
rect 40328 510618 40564 510854
rect 176056 510938 176292 511174
rect 176056 510618 176292 510854
rect 41008 507218 41244 507454
rect 41008 506898 41244 507134
rect 175376 507218 175612 507454
rect 175376 506898 175612 507134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 40328 438938 40564 439174
rect 40328 438618 40564 438854
rect 176056 438938 176292 439174
rect 176056 438618 176292 438854
rect 41008 435218 41244 435454
rect 41008 434898 41244 435134
rect 175376 435218 175612 435454
rect 175376 434898 175612 435134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 40328 402938 40564 403174
rect 40328 402618 40564 402854
rect 176056 402938 176292 403174
rect 176056 402618 176292 402854
rect 41008 399218 41244 399454
rect 41008 398898 41244 399134
rect 175376 399218 175612 399454
rect 175376 398898 175612 399134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 40328 366938 40564 367174
rect 40328 366618 40564 366854
rect 176056 366938 176292 367174
rect 176056 366618 176292 366854
rect 41008 363218 41244 363454
rect 41008 362898 41244 363134
rect 175376 363218 175612 363454
rect 175376 362898 175612 363134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 63866 281258 64102 281494
rect 64186 281258 64422 281494
rect 63866 280938 64102 281174
rect 64186 280938 64422 281174
rect 63866 245258 64102 245494
rect 64186 245258 64422 245494
rect 63866 244938 64102 245174
rect 64186 244938 64422 245174
rect 63866 209258 64102 209494
rect 64186 209258 64422 209494
rect 63866 208938 64102 209174
rect 64186 208938 64422 209174
rect 63866 173258 64102 173494
rect 64186 173258 64422 173494
rect 63866 172938 64102 173174
rect 64186 172938 64422 173174
rect 63866 137258 64102 137494
rect 64186 137258 64422 137494
rect 63866 136938 64102 137174
rect 64186 136938 64422 137174
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 88706 306098 88942 306334
rect 89026 306098 89262 306334
rect 88706 305778 88942 306014
rect 89026 305778 89262 306014
rect 88706 270098 88942 270334
rect 89026 270098 89262 270334
rect 88706 269778 88942 270014
rect 89026 269778 89262 270014
rect 88706 234098 88942 234334
rect 89026 234098 89262 234334
rect 88706 233778 88942 234014
rect 89026 233778 89262 234014
rect 88706 198098 88942 198334
rect 89026 198098 89262 198334
rect 88706 197778 88942 198014
rect 89026 197778 89262 198014
rect 88706 162098 88942 162334
rect 89026 162098 89262 162334
rect 88706 161778 88942 162014
rect 89026 161778 89262 162014
rect 88706 126098 88942 126334
rect 89026 126098 89262 126334
rect 88706 125778 88942 126014
rect 89026 125778 89262 126014
rect 88706 90098 88942 90334
rect 89026 90098 89262 90334
rect 88706 89778 88942 90014
rect 89026 89778 89262 90014
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 92426 309818 92662 310054
rect 92746 309818 92982 310054
rect 92426 309498 92662 309734
rect 92746 309498 92982 309734
rect 92426 273818 92662 274054
rect 92746 273818 92982 274054
rect 92426 273498 92662 273734
rect 92746 273498 92982 273734
rect 92426 237818 92662 238054
rect 92746 237818 92982 238054
rect 92426 237498 92662 237734
rect 92746 237498 92982 237734
rect 92426 201818 92662 202054
rect 92746 201818 92982 202054
rect 92426 201498 92662 201734
rect 92746 201498 92982 201734
rect 92426 165818 92662 166054
rect 92746 165818 92982 166054
rect 92426 165498 92662 165734
rect 92746 165498 92982 165734
rect 92426 129818 92662 130054
rect 92746 129818 92982 130054
rect 92426 129498 92662 129734
rect 92746 129498 92982 129734
rect 92426 93818 92662 94054
rect 92746 93818 92982 94054
rect 92426 93498 92662 93734
rect 92746 93498 92982 93734
rect 92426 57818 92662 58054
rect 92746 57818 92982 58054
rect 92426 57498 92662 57734
rect 92746 57498 92982 57734
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 96146 313538 96382 313774
rect 96466 313538 96702 313774
rect 96146 313218 96382 313454
rect 96466 313218 96702 313454
rect 96146 277538 96382 277774
rect 96466 277538 96702 277774
rect 96146 277218 96382 277454
rect 96466 277218 96702 277454
rect 96146 241538 96382 241774
rect 96466 241538 96702 241774
rect 96146 241218 96382 241454
rect 96466 241218 96702 241454
rect 96146 205538 96382 205774
rect 96466 205538 96702 205774
rect 96146 205218 96382 205454
rect 96466 205218 96702 205454
rect 96146 169538 96382 169774
rect 96466 169538 96702 169774
rect 96146 169218 96382 169454
rect 96466 169218 96702 169454
rect 96146 133538 96382 133774
rect 96466 133538 96702 133774
rect 96146 133218 96382 133454
rect 96466 133218 96702 133454
rect 96146 97538 96382 97774
rect 96466 97538 96702 97774
rect 96146 97218 96382 97454
rect 96466 97218 96702 97454
rect 96146 61538 96382 61774
rect 96466 61538 96702 61774
rect 96146 61218 96382 61454
rect 96466 61218 96702 61454
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 99866 317258 100102 317494
rect 100186 317258 100422 317494
rect 99866 316938 100102 317174
rect 100186 316938 100422 317174
rect 99866 281258 100102 281494
rect 100186 281258 100422 281494
rect 99866 280938 100102 281174
rect 100186 280938 100422 281174
rect 99866 245258 100102 245494
rect 100186 245258 100422 245494
rect 99866 244938 100102 245174
rect 100186 244938 100422 245174
rect 99866 209258 100102 209494
rect 100186 209258 100422 209494
rect 99866 208938 100102 209174
rect 100186 208938 100422 209174
rect 99866 173258 100102 173494
rect 100186 173258 100422 173494
rect 99866 172938 100102 173174
rect 100186 172938 100422 173174
rect 99866 137258 100102 137494
rect 100186 137258 100422 137494
rect 99866 136938 100102 137174
rect 100186 136938 100422 137174
rect 99866 101258 100102 101494
rect 100186 101258 100422 101494
rect 99866 100938 100102 101174
rect 100186 100938 100422 101174
rect 99866 65258 100102 65494
rect 100186 65258 100422 65494
rect 99866 64938 100102 65174
rect 100186 64938 100422 65174
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 124250 183218 124486 183454
rect 124250 182898 124486 183134
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 124250 147218 124486 147454
rect 124250 146898 124486 147134
rect 124706 126098 124942 126334
rect 125026 126098 125262 126334
rect 124706 125778 124942 126014
rect 125026 125778 125262 126014
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 124706 90098 124942 90334
rect 125026 90098 125262 90334
rect 124706 89778 124942 90014
rect 125026 89778 125262 90014
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 128426 165818 128662 166054
rect 128746 165818 128982 166054
rect 128426 165498 128662 165734
rect 128746 165498 128982 165734
rect 128426 129818 128662 130054
rect 128746 129818 128982 130054
rect 128426 129498 128662 129734
rect 128746 129498 128982 129734
rect 128426 93818 128662 94054
rect 128746 93818 128982 94054
rect 128426 93498 128662 93734
rect 128746 93498 128982 93734
rect 128426 57818 128662 58054
rect 128746 57818 128982 58054
rect 128426 57498 128662 57734
rect 128746 57498 128982 57734
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 132146 97538 132382 97774
rect 132466 97538 132702 97774
rect 132146 97218 132382 97454
rect 132466 97218 132702 97454
rect 132146 61538 132382 61774
rect 132466 61538 132702 61774
rect 132146 61218 132382 61454
rect 132466 61218 132702 61454
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 139610 258938 139846 259174
rect 139610 258618 139846 258854
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 139610 222938 139846 223174
rect 139610 222618 139846 222854
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 139610 186938 139846 187174
rect 139610 186618 139846 186854
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 139610 150938 139846 151174
rect 139610 150618 139846 150854
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 139610 114938 139846 115174
rect 139610 114618 139846 114854
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 154970 183218 155206 183454
rect 154970 182898 155206 183134
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 154970 147218 155206 147454
rect 154970 146898 155206 147134
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 170330 258938 170566 259174
rect 170330 258618 170566 258854
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 170330 222938 170566 223174
rect 170330 222618 170566 222854
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 170330 186938 170566 187174
rect 170330 186618 170566 186854
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 170330 150938 170566 151174
rect 170330 150618 170566 150854
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 170330 114938 170566 115174
rect 170330 114618 170566 114854
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 196706 594098 196942 594334
rect 197026 594098 197262 594334
rect 196706 593778 196942 594014
rect 197026 593778 197262 594014
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 200426 597818 200662 598054
rect 200746 597818 200982 598054
rect 200426 597498 200662 597734
rect 200746 597498 200982 597734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 204146 601538 204382 601774
rect 204466 601538 204702 601774
rect 204146 601218 204382 601454
rect 204466 601218 204702 601454
rect 204146 565538 204382 565774
rect 204466 565538 204702 565774
rect 200426 561818 200662 562054
rect 200746 561818 200982 562054
rect 200426 561498 200662 561734
rect 200746 561498 200982 561734
rect 200426 525818 200662 526054
rect 200746 525818 200982 526054
rect 200426 525498 200662 525734
rect 200746 525498 200982 525734
rect 200426 489818 200662 490054
rect 200746 489818 200982 490054
rect 200426 489498 200662 489734
rect 200746 489498 200982 489734
rect 200426 453818 200662 454054
rect 200746 453818 200982 454054
rect 200426 453498 200662 453734
rect 200746 453498 200982 453734
rect 200426 417818 200662 418054
rect 200746 417818 200982 418054
rect 200426 417498 200662 417734
rect 200746 417498 200982 417734
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 204146 565218 204382 565454
rect 204466 565218 204702 565454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 207866 605258 208102 605494
rect 208186 605258 208422 605494
rect 207866 604938 208102 605174
rect 208186 604938 208422 605174
rect 207866 569258 208102 569494
rect 208186 569258 208422 569494
rect 207866 568938 208102 569174
rect 208186 568938 208422 569174
rect 204146 529538 204382 529774
rect 204466 529538 204702 529774
rect 204146 529218 204382 529454
rect 204466 529218 204702 529454
rect 204146 493538 204382 493774
rect 204466 493538 204702 493774
rect 204146 493218 204382 493454
rect 204466 493218 204702 493454
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 204146 421538 204382 421774
rect 204466 421538 204702 421774
rect 204146 421218 204382 421454
rect 204466 421218 204702 421454
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 207866 533258 208102 533494
rect 208186 533258 208422 533494
rect 207866 532938 208102 533174
rect 208186 532938 208422 533174
rect 207866 497258 208102 497494
rect 208186 497258 208422 497494
rect 207866 496938 208102 497174
rect 208186 496938 208422 497174
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 207866 425258 208102 425494
rect 208186 425258 208422 425494
rect 207866 424938 208102 425174
rect 208186 424938 208422 425174
rect 207866 389258 208102 389494
rect 208186 389258 208422 389494
rect 207866 388938 208102 389174
rect 208186 388938 208422 389174
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 220328 654938 220564 655174
rect 220328 654618 220564 654854
rect 356056 654938 356292 655174
rect 356056 654618 356292 654854
rect 221008 651218 221244 651454
rect 221008 650898 221244 651134
rect 355376 651218 355612 651454
rect 355376 650898 355612 651134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 220328 618938 220564 619174
rect 220328 618618 220564 618854
rect 356056 618938 356292 619174
rect 356056 618618 356292 618854
rect 221008 615218 221244 615454
rect 221008 614898 221244 615134
rect 355376 615218 355612 615454
rect 355376 614898 355612 615134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 220328 546938 220564 547174
rect 220328 546618 220564 546854
rect 356056 546938 356292 547174
rect 356056 546618 356292 546854
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 220328 510938 220564 511174
rect 220328 510618 220564 510854
rect 356056 510938 356292 511174
rect 356056 510618 356292 510854
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 220328 438938 220564 439174
rect 220328 438618 220564 438854
rect 356056 438938 356292 439174
rect 356056 438618 356292 438854
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 402938 220564 403174
rect 220328 402618 220564 402854
rect 356056 402938 356292 403174
rect 356056 402618 356292 402854
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 220328 366938 220564 367174
rect 220328 366618 220564 366854
rect 356056 366938 356292 367174
rect 356056 366618 356292 366854
rect 221008 363218 221244 363454
rect 221008 362898 221244 363134
rect 355376 363218 355612 363454
rect 355376 362898 355612 363134
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 240146 349538 240382 349774
rect 240466 349538 240702 349774
rect 240146 349218 240382 349454
rect 240466 349218 240702 349454
rect 240146 313538 240382 313774
rect 240466 313538 240702 313774
rect 240146 313218 240382 313454
rect 240466 313218 240702 313454
rect 243866 353258 244102 353494
rect 244186 353258 244422 353494
rect 243866 352938 244102 353174
rect 244186 352938 244422 353174
rect 243866 317258 244102 317494
rect 244186 317258 244422 317494
rect 243866 316938 244102 317174
rect 244186 316938 244422 317174
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 268706 342098 268942 342334
rect 269026 342098 269262 342334
rect 268706 341778 268942 342014
rect 269026 341778 269262 342014
rect 268706 306098 268942 306334
rect 269026 306098 269262 306334
rect 268706 305778 268942 306014
rect 269026 305778 269262 306014
rect 272426 345818 272662 346054
rect 272746 345818 272982 346054
rect 272426 345498 272662 345734
rect 272746 345498 272982 345734
rect 272426 309818 272662 310054
rect 272746 309818 272982 310054
rect 272426 309498 272662 309734
rect 272746 309498 272982 309734
rect 276146 349538 276382 349774
rect 276466 349538 276702 349774
rect 276146 349218 276382 349454
rect 276466 349218 276702 349454
rect 276146 313538 276382 313774
rect 276466 313538 276702 313774
rect 276146 313218 276382 313454
rect 276466 313218 276702 313454
rect 279866 353258 280102 353494
rect 280186 353258 280422 353494
rect 279866 352938 280102 353174
rect 280186 352938 280422 353174
rect 279866 317258 280102 317494
rect 280186 317258 280422 317494
rect 279866 316938 280102 317174
rect 280186 316938 280422 317174
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 201050 258938 201286 259174
rect 201050 258618 201286 258854
rect 231770 258938 232006 259174
rect 231770 258618 232006 258854
rect 262490 258938 262726 259174
rect 262490 258618 262726 258854
rect 293210 258938 293446 259174
rect 293210 258618 293446 258854
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 216410 255218 216646 255454
rect 216410 254898 216646 255134
rect 247130 255218 247366 255454
rect 247130 254898 247366 255134
rect 277850 255218 278086 255454
rect 277850 254898 278086 255134
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 201050 222938 201286 223174
rect 201050 222618 201286 222854
rect 231770 222938 232006 223174
rect 231770 222618 232006 222854
rect 262490 222938 262726 223174
rect 262490 222618 262726 222854
rect 293210 222938 293446 223174
rect 293210 222618 293446 222854
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 216410 219218 216646 219454
rect 216410 218898 216646 219134
rect 247130 219218 247366 219454
rect 247130 218898 247366 219134
rect 277850 219218 278086 219454
rect 277850 218898 278086 219134
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 201050 186938 201286 187174
rect 201050 186618 201286 186854
rect 231770 186938 232006 187174
rect 231770 186618 232006 186854
rect 262490 186938 262726 187174
rect 262490 186618 262726 186854
rect 293210 186938 293446 187174
rect 293210 186618 293446 186854
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 185690 183218 185926 183454
rect 185690 182898 185926 183134
rect 216410 183218 216646 183454
rect 216410 182898 216646 183134
rect 247130 183218 247366 183454
rect 247130 182898 247366 183134
rect 277850 183218 278086 183454
rect 277850 182898 278086 183134
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 201050 150938 201286 151174
rect 201050 150618 201286 150854
rect 231770 150938 232006 151174
rect 231770 150618 232006 150854
rect 262490 150938 262726 151174
rect 262490 150618 262726 150854
rect 293210 150938 293446 151174
rect 293210 150618 293446 150854
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185690 147218 185926 147454
rect 185690 146898 185926 147134
rect 216410 147218 216646 147454
rect 216410 146898 216646 147134
rect 247130 147218 247366 147454
rect 247130 146898 247366 147134
rect 277850 147218 278086 147454
rect 277850 146898 278086 147134
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 201050 114938 201286 115174
rect 201050 114618 201286 114854
rect 231770 114938 232006 115174
rect 231770 114618 232006 114854
rect 262490 114938 262726 115174
rect 262490 114618 262726 114854
rect 293210 114938 293446 115174
rect 293210 114618 293446 114854
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 216410 111218 216646 111454
rect 216410 110898 216646 111134
rect 247130 111218 247366 111454
rect 247130 110898 247366 111134
rect 277850 111218 278086 111454
rect 277850 110898 278086 111134
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 304706 306098 304942 306334
rect 305026 306098 305262 306334
rect 304706 305778 304942 306014
rect 305026 305778 305262 306014
rect 308426 345818 308662 346054
rect 308746 345818 308982 346054
rect 308426 345498 308662 345734
rect 308746 345498 308982 345734
rect 308426 309818 308662 310054
rect 308746 309818 308982 310054
rect 308426 309498 308662 309734
rect 308746 309498 308982 309734
rect 312146 349538 312382 349774
rect 312466 349538 312702 349774
rect 312146 349218 312382 349454
rect 312466 349218 312702 349454
rect 312146 313538 312382 313774
rect 312466 313538 312702 313774
rect 312146 313218 312382 313454
rect 312466 313218 312702 313454
rect 304706 270098 304942 270334
rect 305026 270098 305262 270334
rect 304706 269778 304942 270014
rect 305026 269778 305262 270014
rect 312146 277538 312382 277774
rect 312466 277538 312702 277774
rect 312146 277218 312382 277454
rect 312466 277218 312702 277454
rect 308570 255218 308806 255454
rect 308570 254898 308806 255134
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 308570 219218 308806 219454
rect 308570 218898 308806 219134
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 308570 183218 308806 183454
rect 308570 182898 308806 183134
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 308570 147218 308806 147454
rect 308570 146898 308806 147134
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 308570 111218 308806 111454
rect 308570 110898 308806 111134
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 353258 316102 353494
rect 316186 353258 316422 353494
rect 315866 352938 316102 353174
rect 316186 352938 316422 353174
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 342098 340942 342334
rect 341026 342098 341262 342334
rect 340706 341778 340942 342014
rect 341026 341778 341262 342014
rect 340706 306098 340942 306334
rect 341026 306098 341262 306334
rect 340706 305778 340942 306014
rect 341026 305778 341262 306014
rect 340706 270098 340942 270334
rect 341026 270098 341262 270334
rect 340706 269778 340942 270014
rect 341026 269778 341262 270014
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 340706 90098 340942 90334
rect 341026 90098 341262 90334
rect 340706 89778 340942 90014
rect 341026 89778 341262 90014
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 345818 344662 346054
rect 344746 345818 344982 346054
rect 344426 345498 344662 345734
rect 344746 345498 344982 345734
rect 344426 309818 344662 310054
rect 344746 309818 344982 310054
rect 344426 309498 344662 309734
rect 344746 309498 344982 309734
rect 344426 273818 344662 274054
rect 344746 273818 344982 274054
rect 344426 273498 344662 273734
rect 344746 273498 344982 273734
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 349538 348382 349774
rect 348466 349538 348702 349774
rect 348146 349218 348382 349454
rect 348466 349218 348702 349454
rect 348146 313538 348382 313774
rect 348466 313538 348702 313774
rect 348146 313218 348382 313454
rect 348466 313218 348702 313454
rect 348146 277538 348382 277774
rect 348466 277538 348702 277774
rect 348146 277218 348382 277454
rect 348466 277218 348702 277454
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 353258 352102 353494
rect 352186 353258 352422 353494
rect 351866 352938 352102 353174
rect 352186 352938 352422 353174
rect 351866 317258 352102 317494
rect 352186 317258 352422 317494
rect 351866 316938 352102 317174
rect 352186 316938 352422 317174
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 351866 281258 352102 281494
rect 352186 281258 352422 281494
rect 351866 280938 352102 281174
rect 352186 280938 352422 281174
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 364250 219218 364486 219454
rect 364250 218898 364486 219134
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 364250 183218 364486 183454
rect 364250 182898 364486 183134
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 364250 147218 364486 147454
rect 364250 146898 364486 147134
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 364250 111218 364486 111454
rect 364250 110898 364486 111134
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 364250 75218 364486 75454
rect 364250 74898 364486 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 379610 222938 379846 223174
rect 379610 222618 379846 222854
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 379610 186938 379846 187174
rect 379610 186618 379846 186854
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 379610 150938 379846 151174
rect 379610 150618 379846 150854
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 379610 114938 379846 115174
rect 379610 114618 379846 114854
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 379610 78938 379846 79174
rect 379610 78618 379846 78854
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 400328 654938 400564 655174
rect 400328 654618 400564 654854
rect 536056 654938 536292 655174
rect 536056 654618 536292 654854
rect 401008 651218 401244 651454
rect 401008 650898 401244 651134
rect 535376 651218 535612 651454
rect 535376 650898 535612 651134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 400328 618938 400564 619174
rect 400328 618618 400564 618854
rect 536056 618938 536292 619174
rect 536056 618618 536292 618854
rect 401008 615218 401244 615454
rect 401008 614898 401244 615134
rect 535376 615218 535612 615454
rect 535376 614898 535612 615134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 400328 546938 400564 547174
rect 400328 546618 400564 546854
rect 536056 546938 536292 547174
rect 536056 546618 536292 546854
rect 401008 543218 401244 543454
rect 401008 542898 401244 543134
rect 535376 543218 535612 543454
rect 535376 542898 535612 543134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 400328 510938 400564 511174
rect 400328 510618 400564 510854
rect 536056 510938 536292 511174
rect 536056 510618 536292 510854
rect 401008 507218 401244 507454
rect 401008 506898 401244 507134
rect 535376 507218 535612 507454
rect 535376 506898 535612 507134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 400328 438938 400564 439174
rect 400328 438618 400564 438854
rect 536056 438938 536292 439174
rect 536056 438618 536292 438854
rect 401008 435218 401244 435454
rect 401008 434898 401244 435134
rect 535376 435218 535612 435454
rect 535376 434898 535612 435134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 400328 402938 400564 403174
rect 400328 402618 400564 402854
rect 536056 402938 536292 403174
rect 536056 402618 536292 402854
rect 401008 399218 401244 399454
rect 401008 398898 401244 399134
rect 535376 399218 535612 399454
rect 535376 398898 535612 399134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 400328 366938 400564 367174
rect 400328 366618 400564 366854
rect 536056 366938 536292 367174
rect 536056 366618 536292 366854
rect 401008 363218 401244 363454
rect 401008 362898 401244 363134
rect 535376 363218 535612 363454
rect 535376 362898 535612 363134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 394970 219218 395206 219454
rect 394970 218898 395206 219134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 394970 183218 395206 183454
rect 394970 182898 395206 183134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 394970 147218 395206 147454
rect 394970 146898 395206 147134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 394970 111218 395206 111454
rect 394970 110898 395206 111134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 394970 75218 395206 75454
rect 394970 74898 395206 75134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 484706 234098 484942 234334
rect 485026 234098 485262 234334
rect 484706 233778 484942 234014
rect 485026 233778 485262 234014
rect 488426 345818 488662 346054
rect 488746 345818 488982 346054
rect 488426 345498 488662 345734
rect 488746 345498 488982 345734
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 488426 237818 488662 238054
rect 488746 237818 488982 238054
rect 488426 237498 488662 237734
rect 488746 237498 488982 237734
rect 492146 349538 492382 349774
rect 492466 349538 492702 349774
rect 492146 349218 492382 349454
rect 492466 349218 492702 349454
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 492146 241538 492382 241774
rect 492466 241538 492702 241774
rect 492146 241218 492382 241454
rect 492466 241218 492702 241454
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 410330 222938 410566 223174
rect 410330 222618 410566 222854
rect 441050 222938 441286 223174
rect 441050 222618 441286 222854
rect 471770 222938 472006 223174
rect 471770 222618 472006 222854
rect 425690 219218 425926 219454
rect 425690 218898 425926 219134
rect 456410 219218 456646 219454
rect 456410 218898 456646 219134
rect 487130 219218 487366 219454
rect 487130 218898 487366 219134
rect 492146 205538 492382 205774
rect 492466 205538 492702 205774
rect 492146 205218 492382 205454
rect 492466 205218 492702 205454
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 410330 186938 410566 187174
rect 410330 186618 410566 186854
rect 441050 186938 441286 187174
rect 441050 186618 441286 186854
rect 471770 186938 472006 187174
rect 471770 186618 472006 186854
rect 425690 183218 425926 183454
rect 425690 182898 425926 183134
rect 456410 183218 456646 183454
rect 456410 182898 456646 183134
rect 487130 183218 487366 183454
rect 487130 182898 487366 183134
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 410330 150938 410566 151174
rect 410330 150618 410566 150854
rect 441050 150938 441286 151174
rect 441050 150618 441286 150854
rect 471770 150938 472006 151174
rect 471770 150618 472006 150854
rect 425690 147218 425926 147454
rect 425690 146898 425926 147134
rect 456410 147218 456646 147454
rect 456410 146898 456646 147134
rect 487130 147218 487366 147454
rect 487130 146898 487366 147134
rect 492146 133538 492382 133774
rect 492466 133538 492702 133774
rect 492146 133218 492382 133454
rect 492466 133218 492702 133454
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 410330 114938 410566 115174
rect 410330 114618 410566 114854
rect 441050 114938 441286 115174
rect 441050 114618 441286 114854
rect 471770 114938 472006 115174
rect 471770 114618 472006 114854
rect 425690 111218 425926 111454
rect 425690 110898 425926 111134
rect 456410 111218 456646 111454
rect 456410 110898 456646 111134
rect 487130 111218 487366 111454
rect 487130 110898 487366 111134
rect 492146 97538 492382 97774
rect 492466 97538 492702 97774
rect 492146 97218 492382 97454
rect 492466 97218 492702 97454
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 410330 78938 410566 79174
rect 410330 78618 410566 78854
rect 441050 78938 441286 79174
rect 441050 78618 441286 78854
rect 471770 78938 472006 79174
rect 471770 78618 472006 78854
rect 425690 75218 425926 75454
rect 425690 74898 425926 75134
rect 456410 75218 456646 75454
rect 456410 74898 456646 75134
rect 487130 75218 487366 75454
rect 487130 74898 487366 75134
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 495866 245258 496102 245494
rect 496186 245258 496422 245494
rect 495866 244938 496102 245174
rect 496186 244938 496422 245174
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 502490 222938 502726 223174
rect 502490 222618 502726 222854
rect 495866 209258 496102 209494
rect 496186 209258 496422 209494
rect 495866 208938 496102 209174
rect 496186 208938 496422 209174
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 502490 186938 502726 187174
rect 502490 186618 502726 186854
rect 495866 173258 496102 173494
rect 496186 173258 496422 173494
rect 495866 172938 496102 173174
rect 496186 172938 496422 173174
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 502490 150938 502726 151174
rect 502490 150618 502726 150854
rect 495866 137258 496102 137494
rect 496186 137258 496422 137494
rect 495866 136938 496102 137174
rect 496186 136938 496422 137174
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 502490 114938 502726 115174
rect 502490 114618 502726 114854
rect 495866 101258 496102 101494
rect 496186 101258 496422 101494
rect 495866 100938 496102 101174
rect 496186 100938 496422 101174
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 502490 78938 502726 79174
rect 502490 78618 502726 78854
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 517850 219218 518086 219454
rect 517850 218898 518086 219134
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 517850 183218 518086 183454
rect 517850 182898 518086 183134
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 517850 147218 518086 147454
rect 517850 146898 518086 147134
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 520706 126098 520942 126334
rect 521026 126098 521262 126334
rect 520706 125778 520942 126014
rect 521026 125778 521262 126014
rect 517850 111218 518086 111454
rect 517850 110898 518086 111134
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 520706 90098 520942 90334
rect 521026 90098 521262 90334
rect 520706 89778 520942 90014
rect 521026 89778 521262 90014
rect 517850 75218 518086 75454
rect 517850 74898 518086 75134
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 524426 129818 524662 130054
rect 524746 129818 524982 130054
rect 524426 129498 524662 129734
rect 524746 129498 524982 129734
rect 524426 93818 524662 94054
rect 524746 93818 524982 94054
rect 524426 93498 524662 93734
rect 524746 93498 524982 93734
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 528146 133538 528382 133774
rect 528466 133538 528702 133774
rect 528146 133218 528382 133454
rect 528466 133218 528702 133454
rect 528146 97538 528382 97774
rect 528466 97538 528702 97774
rect 528146 97218 528382 97454
rect 528466 97218 528702 97454
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 533210 222938 533446 223174
rect 533210 222618 533446 222854
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 533210 186938 533446 187174
rect 533210 186618 533446 186854
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 533210 150938 533446 151174
rect 533210 150618 533446 150854
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 533210 114938 533446 115174
rect 533210 114618 533446 114854
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 533210 78938 533446 79174
rect 533210 78618 533446 78854
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 40328 655174
rect 40564 654938 176056 655174
rect 176292 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 220328 655174
rect 220564 654938 356056 655174
rect 356292 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 400328 655174
rect 400564 654938 536056 655174
rect 536292 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 40328 654854
rect 40564 654618 176056 654854
rect 176292 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 220328 654854
rect 220564 654618 356056 654854
rect 356292 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 400328 654854
rect 400564 654618 536056 654854
rect 536292 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 41008 651454
rect 41244 651218 175376 651454
rect 175612 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 221008 651454
rect 221244 651218 355376 651454
rect 355612 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 401008 651454
rect 401244 651218 535376 651454
rect 535612 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 41008 651134
rect 41244 650898 175376 651134
rect 175612 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 221008 651134
rect 221244 650898 355376 651134
rect 355612 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 401008 651134
rect 401244 650898 535376 651134
rect 535612 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 40328 619174
rect 40564 618938 176056 619174
rect 176292 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 220328 619174
rect 220564 618938 356056 619174
rect 356292 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 400328 619174
rect 400564 618938 536056 619174
rect 536292 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 40328 618854
rect 40564 618618 176056 618854
rect 176292 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 220328 618854
rect 220564 618618 356056 618854
rect 356292 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 400328 618854
rect 400564 618618 536056 618854
rect 536292 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 41008 615454
rect 41244 615218 175376 615454
rect 175612 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 221008 615454
rect 221244 615218 355376 615454
rect 355612 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 401008 615454
rect 401244 615218 535376 615454
rect 535612 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 41008 615134
rect 41244 614898 175376 615134
rect 175612 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 221008 615134
rect 221244 614898 355376 615134
rect 355612 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 401008 615134
rect 401244 614898 535376 615134
rect 535612 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 40328 547174
rect 40564 546938 176056 547174
rect 176292 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 220328 547174
rect 220564 546938 356056 547174
rect 356292 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 400328 547174
rect 400564 546938 536056 547174
rect 536292 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 40328 546854
rect 40564 546618 176056 546854
rect 176292 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 220328 546854
rect 220564 546618 356056 546854
rect 356292 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 400328 546854
rect 400564 546618 536056 546854
rect 536292 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 41008 543454
rect 41244 543218 175376 543454
rect 175612 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 401008 543454
rect 401244 543218 535376 543454
rect 535612 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 41008 543134
rect 41244 542898 175376 543134
rect 175612 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 401008 543134
rect 401244 542898 535376 543134
rect 535612 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 40328 511174
rect 40564 510938 176056 511174
rect 176292 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 220328 511174
rect 220564 510938 356056 511174
rect 356292 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 400328 511174
rect 400564 510938 536056 511174
rect 536292 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 40328 510854
rect 40564 510618 176056 510854
rect 176292 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 220328 510854
rect 220564 510618 356056 510854
rect 356292 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 400328 510854
rect 400564 510618 536056 510854
rect 536292 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 41008 507454
rect 41244 507218 175376 507454
rect 175612 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 401008 507454
rect 401244 507218 535376 507454
rect 535612 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 41008 507134
rect 41244 506898 175376 507134
rect 175612 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 401008 507134
rect 401244 506898 535376 507134
rect 535612 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 40328 439174
rect 40564 438938 176056 439174
rect 176292 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 220328 439174
rect 220564 438938 356056 439174
rect 356292 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 400328 439174
rect 400564 438938 536056 439174
rect 536292 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 40328 438854
rect 40564 438618 176056 438854
rect 176292 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 220328 438854
rect 220564 438618 356056 438854
rect 356292 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 400328 438854
rect 400564 438618 536056 438854
rect 536292 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 41008 435454
rect 41244 435218 175376 435454
rect 175612 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 401008 435454
rect 401244 435218 535376 435454
rect 535612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 41008 435134
rect 41244 434898 175376 435134
rect 175612 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 401008 435134
rect 401244 434898 535376 435134
rect 535612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 40328 403174
rect 40564 402938 176056 403174
rect 176292 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 220328 403174
rect 220564 402938 356056 403174
rect 356292 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 400328 403174
rect 400564 402938 536056 403174
rect 536292 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 40328 402854
rect 40564 402618 176056 402854
rect 176292 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 220328 402854
rect 220564 402618 356056 402854
rect 356292 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 400328 402854
rect 400564 402618 536056 402854
rect 536292 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 41008 399454
rect 41244 399218 175376 399454
rect 175612 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 401008 399454
rect 401244 399218 535376 399454
rect 535612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 41008 399134
rect 41244 398898 175376 399134
rect 175612 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 401008 399134
rect 401244 398898 535376 399134
rect 535612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 40328 367174
rect 40564 366938 176056 367174
rect 176292 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 220328 367174
rect 220564 366938 356056 367174
rect 356292 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 400328 367174
rect 400564 366938 536056 367174
rect 536292 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 40328 366854
rect 40564 366618 176056 366854
rect 176292 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 220328 366854
rect 220564 366618 356056 366854
rect 356292 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 400328 366854
rect 400564 366618 536056 366854
rect 536292 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 41008 363454
rect 41244 363218 175376 363454
rect 175612 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 221008 363454
rect 221244 363218 355376 363454
rect 355612 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 401008 363454
rect 401244 363218 535376 363454
rect 535612 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 41008 363134
rect 41244 362898 175376 363134
rect 175612 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 221008 363134
rect 221244 362898 355376 363134
rect 355612 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 401008 363134
rect 401244 362898 535376 363134
rect 535612 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 276146 313774
rect 276382 313538 276466 313774
rect 276702 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 276146 313454
rect 276382 313218 276466 313454
rect 276702 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 272426 310054
rect 272662 309818 272746 310054
rect 272982 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 272426 309734
rect 272662 309498 272746 309734
rect 272982 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 268706 306334
rect 268942 306098 269026 306334
rect 269262 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 268706 306014
rect 268942 305778 269026 306014
rect 269262 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 139610 259174
rect 139846 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 170330 259174
rect 170566 258938 201050 259174
rect 201286 258938 231770 259174
rect 232006 258938 262490 259174
rect 262726 258938 293210 259174
rect 293446 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 139610 258854
rect 139846 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 170330 258854
rect 170566 258618 201050 258854
rect 201286 258618 231770 258854
rect 232006 258618 262490 258854
rect 262726 258618 293210 258854
rect 293446 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 154970 255454
rect 155206 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 185690 255454
rect 185926 255218 216410 255454
rect 216646 255218 247130 255454
rect 247366 255218 277850 255454
rect 278086 255218 308570 255454
rect 308806 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 154970 255134
rect 155206 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 185690 255134
rect 185926 254898 216410 255134
rect 216646 254898 247130 255134
rect 247366 254898 277850 255134
rect 278086 254898 308570 255134
rect 308806 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 139610 223174
rect 139846 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 170330 223174
rect 170566 222938 201050 223174
rect 201286 222938 231770 223174
rect 232006 222938 262490 223174
rect 262726 222938 293210 223174
rect 293446 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 379610 223174
rect 379846 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 410330 223174
rect 410566 222938 441050 223174
rect 441286 222938 471770 223174
rect 472006 222938 502490 223174
rect 502726 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 533210 223174
rect 533446 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 139610 222854
rect 139846 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 170330 222854
rect 170566 222618 201050 222854
rect 201286 222618 231770 222854
rect 232006 222618 262490 222854
rect 262726 222618 293210 222854
rect 293446 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 379610 222854
rect 379846 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 410330 222854
rect 410566 222618 441050 222854
rect 441286 222618 471770 222854
rect 472006 222618 502490 222854
rect 502726 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 533210 222854
rect 533446 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 154970 219454
rect 155206 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 185690 219454
rect 185926 219218 216410 219454
rect 216646 219218 247130 219454
rect 247366 219218 277850 219454
rect 278086 219218 308570 219454
rect 308806 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 364250 219454
rect 364486 219218 394970 219454
rect 395206 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 425690 219454
rect 425926 219218 456410 219454
rect 456646 219218 487130 219454
rect 487366 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 517850 219454
rect 518086 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 154970 219134
rect 155206 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 185690 219134
rect 185926 218898 216410 219134
rect 216646 218898 247130 219134
rect 247366 218898 277850 219134
rect 278086 218898 308570 219134
rect 308806 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 364250 219134
rect 364486 218898 394970 219134
rect 395206 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 425690 219134
rect 425926 218898 456410 219134
rect 456646 218898 487130 219134
rect 487366 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 517850 219134
rect 518086 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 139610 187174
rect 139846 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 170330 187174
rect 170566 186938 201050 187174
rect 201286 186938 231770 187174
rect 232006 186938 262490 187174
rect 262726 186938 293210 187174
rect 293446 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 379610 187174
rect 379846 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 410330 187174
rect 410566 186938 441050 187174
rect 441286 186938 471770 187174
rect 472006 186938 502490 187174
rect 502726 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 533210 187174
rect 533446 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 139610 186854
rect 139846 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 170330 186854
rect 170566 186618 201050 186854
rect 201286 186618 231770 186854
rect 232006 186618 262490 186854
rect 262726 186618 293210 186854
rect 293446 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 379610 186854
rect 379846 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 410330 186854
rect 410566 186618 441050 186854
rect 441286 186618 471770 186854
rect 472006 186618 502490 186854
rect 502726 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 533210 186854
rect 533446 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 124250 183454
rect 124486 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 154970 183454
rect 155206 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 185690 183454
rect 185926 183218 216410 183454
rect 216646 183218 247130 183454
rect 247366 183218 277850 183454
rect 278086 183218 308570 183454
rect 308806 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 364250 183454
rect 364486 183218 394970 183454
rect 395206 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 425690 183454
rect 425926 183218 456410 183454
rect 456646 183218 487130 183454
rect 487366 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 517850 183454
rect 518086 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 124250 183134
rect 124486 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 154970 183134
rect 155206 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 185690 183134
rect 185926 182898 216410 183134
rect 216646 182898 247130 183134
rect 247366 182898 277850 183134
rect 278086 182898 308570 183134
rect 308806 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 364250 183134
rect 364486 182898 394970 183134
rect 395206 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 425690 183134
rect 425926 182898 456410 183134
rect 456646 182898 487130 183134
rect 487366 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 517850 183134
rect 518086 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 139610 151174
rect 139846 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 170330 151174
rect 170566 150938 201050 151174
rect 201286 150938 231770 151174
rect 232006 150938 262490 151174
rect 262726 150938 293210 151174
rect 293446 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 379610 151174
rect 379846 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 410330 151174
rect 410566 150938 441050 151174
rect 441286 150938 471770 151174
rect 472006 150938 502490 151174
rect 502726 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 533210 151174
rect 533446 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 139610 150854
rect 139846 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 170330 150854
rect 170566 150618 201050 150854
rect 201286 150618 231770 150854
rect 232006 150618 262490 150854
rect 262726 150618 293210 150854
rect 293446 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 379610 150854
rect 379846 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 410330 150854
rect 410566 150618 441050 150854
rect 441286 150618 471770 150854
rect 472006 150618 502490 150854
rect 502726 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 533210 150854
rect 533446 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 124250 147454
rect 124486 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 154970 147454
rect 155206 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 185690 147454
rect 185926 147218 216410 147454
rect 216646 147218 247130 147454
rect 247366 147218 277850 147454
rect 278086 147218 308570 147454
rect 308806 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 364250 147454
rect 364486 147218 394970 147454
rect 395206 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 425690 147454
rect 425926 147218 456410 147454
rect 456646 147218 487130 147454
rect 487366 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 517850 147454
rect 518086 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 124250 147134
rect 124486 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 154970 147134
rect 155206 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 185690 147134
rect 185926 146898 216410 147134
rect 216646 146898 247130 147134
rect 247366 146898 277850 147134
rect 278086 146898 308570 147134
rect 308806 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 364250 147134
rect 364486 146898 394970 147134
rect 395206 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 425690 147134
rect 425926 146898 456410 147134
rect 456646 146898 487130 147134
rect 487366 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 517850 147134
rect 518086 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 139610 115174
rect 139846 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 170330 115174
rect 170566 114938 201050 115174
rect 201286 114938 231770 115174
rect 232006 114938 262490 115174
rect 262726 114938 293210 115174
rect 293446 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 379610 115174
rect 379846 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 410330 115174
rect 410566 114938 441050 115174
rect 441286 114938 471770 115174
rect 472006 114938 502490 115174
rect 502726 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 533210 115174
rect 533446 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 139610 114854
rect 139846 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 170330 114854
rect 170566 114618 201050 114854
rect 201286 114618 231770 114854
rect 232006 114618 262490 114854
rect 262726 114618 293210 114854
rect 293446 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 379610 114854
rect 379846 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 410330 114854
rect 410566 114618 441050 114854
rect 441286 114618 471770 114854
rect 472006 114618 502490 114854
rect 502726 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 533210 114854
rect 533446 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 154970 111454
rect 155206 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 185690 111454
rect 185926 111218 216410 111454
rect 216646 111218 247130 111454
rect 247366 111218 277850 111454
rect 278086 111218 308570 111454
rect 308806 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 364250 111454
rect 364486 111218 394970 111454
rect 395206 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 425690 111454
rect 425926 111218 456410 111454
rect 456646 111218 487130 111454
rect 487366 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 517850 111454
rect 518086 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 154970 111134
rect 155206 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 185690 111134
rect 185926 110898 216410 111134
rect 216646 110898 247130 111134
rect 247366 110898 277850 111134
rect 278086 110898 308570 111134
rect 308806 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 364250 111134
rect 364486 110898 394970 111134
rect 395206 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 425690 111134
rect 425926 110898 456410 111134
rect 456646 110898 487130 111134
rect 487366 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 517850 111134
rect 518086 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 379610 79174
rect 379846 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 410330 79174
rect 410566 78938 441050 79174
rect 441286 78938 471770 79174
rect 472006 78938 502490 79174
rect 502726 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 533210 79174
rect 533446 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 379610 78854
rect 379846 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 410330 78854
rect 410566 78618 441050 78854
rect 441286 78618 471770 78854
rect 472006 78618 502490 78854
rect 502726 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 533210 78854
rect 533446 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 364250 75454
rect 364486 75218 394970 75454
rect 395206 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 425690 75454
rect 425926 75218 456410 75454
rect 456646 75218 487130 75454
rect 487366 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 517850 75454
rect 518086 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 364250 75134
rect 364486 74898 394970 75134
rect 395206 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 425690 75134
rect 425926 74898 456410 75134
rect 456646 74898 487130 75134
rect 487366 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 517850 75134
rect 518086 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use io_interface  IO_interface
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 198850 200000
use sky130_sram_2kbyte_1rw1r_32x512_8  data_memory
timestamp 0
transform 1 0 40000 0 1 360000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory0
timestamp 0
transform 1 0 40000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory1
timestamp 0
transform 1 0 40000 0 1 600000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory2
timestamp 0
transform 1 0 220000 0 1 360000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory3
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory4
timestamp 0
transform 1 0 220000 0 1 600000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory5
timestamp 0
transform 1 0 400000 0 1 360000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory6
timestamp 0
transform 1 0 400000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory7
timestamp 0
transform 1 0 400000 0 1 600000
box 0 0 136620 83308
use processor  uP
timestamp 0
transform 1 0 360000 0 1 50000
box 1066 0 178886 180000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 685244 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 685244 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 685244 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 357940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 685244 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 79743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 281537 218414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 685244 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 79743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 281537 254414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 685244 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 79743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 281537 290414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 685244 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 357940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 685244 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 685244 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 51375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 228961 434414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 685244 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 51375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 228961 470414 358064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 685244 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 357940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 685244 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 685244 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 357940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 685244 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 685244 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 685244 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 79743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 281537 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 79743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 281537 225854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 685244 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 79743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 281537 261854 357940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 685244 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 685244 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 685244 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 51375 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 228961 405854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 685244 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 50068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 229452 441854 357940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 685244 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 51375 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 228961 477854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 685244 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 358064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 685244 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 357940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 79743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 281537 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 79743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 281537 233294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 79743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 281537 269294 357940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 51375 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 228961 413294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 51375 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 228961 449294 357940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 51375 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 228961 485294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 358064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 357940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 357940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 358064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 358064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 79743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 281537 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 79743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 281537 240734 357940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 79743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 281537 276734 357940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 358064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 358064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 51375 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 228961 420734 357940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 50068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 229452 456734 357940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 358064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 358064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 357940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 79743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 281537 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 79743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 281537 237014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 79743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 281537 273014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 80068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 279580 309014 357940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 51375 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 228961 417014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 51375 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 228961 453014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 51375 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 228961 489014 357940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 358064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 357940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 358064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 357940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 358064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 79743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 281537 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 79743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 281537 244454 357940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 79743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 281537 280454 358064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 357940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 358064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 51375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 228961 424454 357940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 51375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 228961 460454 358064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 357940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 358064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 358064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 685244 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 357940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 685244 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 357940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 685244 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 358064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 685244 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 79743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 281537 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 79743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 281537 222134 358064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 685244 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 79743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 281537 258134 357940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 685244 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 79743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 281537 294134 357940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 685244 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 358064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 685244 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 358064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 685244 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 51375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 228961 438134 357940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 685244 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 51375 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 228961 474134 357940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 685244 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 358064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 685244 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 358064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 685244 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 357940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 685244 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 357940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 685244 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 358064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 685244 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 79743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 281537 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 79743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 281537 229574 358064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 685244 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 79743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 281537 265574 357940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 685244 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 357940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 685244 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 358064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 685244 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 51375 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 228961 409574 358064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 685244 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 51375 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 228961 445574 357940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 685244 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 51375 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 228961 481574 357940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 685244 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 358064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 685244 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 535494 651336 535494 651336 0 vccd1
rlabel via4 513704 226776 513704 226776 0 vccd2
rlabel via4 521144 198216 521144 198216 0 vdda1
rlabel via4 528584 205656 528584 205656 0 vdda2
rlabel via4 524864 201936 524864 201936 0 vssa1
rlabel via4 532304 209376 532304 209376 0 vssa2
rlabel via4 536174 655056 536174 655056 0 vssd1
rlabel via4 517424 194496 517424 194496 0 vssd2
rlabel via1 314134 80597 314134 80597 0 Serial_input
rlabel metal2 315514 79271 315514 79271 0 Serial_output
rlabel metal3 40020 368360 40020 368360 0 clk
rlabel metal3 56281 357340 56281 357340 0 data_mem_addr\[0\]
rlabel metal3 57891 357204 57891 357204 0 data_mem_addr\[1\]
rlabel metal3 39353 387804 39353 387804 0 data_mem_addr\[2\]
rlabel metal3 39399 389436 39399 389436 0 data_mem_addr\[3\]
rlabel metal3 39491 390660 39491 390660 0 data_mem_addr\[4\]
rlabel metal3 39445 392292 39445 392292 0 data_mem_addr\[5\]
rlabel metal3 39537 393516 39537 393516 0 data_mem_addr\[6\]
rlabel metal3 39261 395420 39261 395420 0 data_mem_addr\[7\]
rlabel metal3 39215 367540 39215 367540 0 data_mem_csb
rlabel metal2 192158 279956 192158 279956 0 data_read_data\[0\]
rlabel metal1 148212 349826 148212 349826 0 data_read_data\[10\]
rlabel metal3 96255 357340 96255 357340 0 data_read_data\[11\]
rlabel metal3 98923 357340 98923 357340 0 data_read_data\[12\]
rlabel metal3 101499 357340 101499 357340 0 data_read_data\[13\]
rlabel metal4 103316 357748 103316 357748 0 data_read_data\[14\]
rlabel metal1 156722 307122 156722 307122 0 data_read_data\[15\]
rlabel metal2 193630 279956 193630 279956 0 data_read_data\[1\]
rlabel metal2 195102 279956 195102 279956 0 data_read_data\[2\]
rlabel metal2 77234 356337 77234 356337 0 data_read_data\[3\]
rlabel metal3 78545 357340 78545 357340 0 data_read_data\[4\]
rlabel metal3 81213 357340 81213 357340 0 data_read_data\[5\]
rlabel metal3 83881 356660 83881 356660 0 data_read_data\[6\]
rlabel metal1 144118 293318 144118 293318 0 data_read_data\[7\]
rlabel metal1 145176 313990 145176 313990 0 data_read_data\[8\]
rlabel metal1 146924 315350 146924 315350 0 data_read_data\[9\]
rlabel metal3 58765 357340 58765 357340 0 data_wmask\[0\]
rlabel metal1 61732 356626 61732 356626 0 data_wmask\[1\]
rlabel metal3 61019 358156 61019 358156 0 data_wmask\[2\]
rlabel metal3 61985 357340 61985 357340 0 data_wmask\[3\]
rlabel metal3 63319 357340 63319 357340 0 data_write_data\[0\]
rlabel metal3 75233 357340 75233 357340 0 data_write_data\[10\]
rlabel metal3 76475 357204 76475 357204 0 data_write_data\[11\]
rlabel metal3 76521 357340 76521 357340 0 data_write_data\[12\]
rlabel metal3 78407 357204 78407 357204 0 data_write_data\[13\]
rlabel metal3 79787 357340 79787 357340 0 data_write_data\[14\]
rlabel metal3 80983 357204 80983 357204 0 data_write_data\[15\]
rlabel metal2 64354 357119 64354 357119 0 data_write_data\[1\]
rlabel metal4 64676 357748 64676 357748 0 data_write_data\[2\]
rlabel metal2 197310 279956 197310 279956 0 data_write_data\[3\]
rlabel metal2 198414 279956 198414 279956 0 data_write_data\[4\]
rlabel metal2 199518 279956 199518 279956 0 data_write_data\[5\]
rlabel metal1 135470 329154 135470 329154 0 data_write_data\[6\]
rlabel metal1 136804 296106 136804 296106 0 data_write_data\[7\]
rlabel metal3 72749 357340 72749 357340 0 data_write_data\[8\]
rlabel metal2 74106 356677 74106 356677 0 data_write_data\[9\]
rlabel metal3 39307 369852 39307 369852 0 dataw_enb
rlabel metal2 312754 79339 312754 79339 0 hlt
rlabel metal2 55430 596445 55430 596445 0 instr_mem_addr_9bit\[0\]
rlabel metal2 39928 485044 39928 485044 0 instr_mem_addr_9bit\[1\]
rlabel metal3 38042 507892 38042 507892 0 instr_mem_addr_9bit\[2\]
rlabel metal3 40020 509930 40020 509930 0 instr_mem_addr_9bit\[3\]
rlabel metal3 40020 511018 40020 511018 0 instr_mem_addr_9bit\[4\]
rlabel metal3 40020 513088 40020 513088 0 instr_mem_addr_9bit\[5\]
rlabel metal3 40020 513904 40020 513904 0 instr_mem_addr_9bit\[6\]
rlabel metal1 38134 585174 38134 585174 0 instr_mem_addr_9bit\[7\]
rlabel metal3 38939 636276 38939 636276 0 instr_mem_addr_9bit\[8\]
rlabel metal3 39468 487492 39468 487492 0 instr_mem_csb\[0\]
rlabel metal3 39376 607444 39376 607444 0 instr_mem_csb\[1\]
rlabel metal2 217442 361641 217442 361641 0 instr_mem_csb\[2\]
rlabel metal1 222410 353974 222410 353974 0 instr_mem_csb\[3\]
rlabel metal2 221966 279956 221966 279956 0 instr_mem_csb\[4\]
rlabel metal2 217550 279956 217550 279956 0 instr_mem_csb\[5\]
rlabel metal2 213134 279956 213134 279956 0 instr_mem_csb\[6\]
rlabel metal3 283337 294508 283337 294508 0 instr_mem_csb\[7\]
rlabel metal1 138782 445026 138782 445026 0 instr_read_data0\[0\]
rlabel via3 216867 369852 216867 369852 0 instr_read_data0\[10\]
rlabel metal3 96347 476204 96347 476204 0 instr_read_data0\[11\]
rlabel metal3 98923 476204 98923 476204 0 instr_read_data0\[12\]
rlabel metal3 101499 476204 101499 476204 0 instr_read_data0\[13\]
rlabel metal4 103316 478176 103316 478176 0 instr_read_data0\[14\]
rlabel metal2 215050 365177 215050 365177 0 instr_read_data0\[15\]
rlabel metal4 214636 366452 214636 366452 0 instr_read_data0\[16\]
rlabel metal4 214820 366452 214820 366452 0 instr_read_data0\[17\]
rlabel metal3 113965 476204 113965 476204 0 instr_read_data0\[18\]
rlabel metal3 116633 476204 116633 476204 0 instr_read_data0\[19\]
rlabel metal2 213410 279956 213410 279956 0 instr_read_data0\[1\]
rlabel via3 118611 476204 118611 476204 0 instr_read_data0\[20\]
rlabel metal3 121187 476204 121187 476204 0 instr_read_data0\[21\]
rlabel metal2 212290 368390 212290 368390 0 instr_read_data0\[22\]
rlabel metal2 212106 367982 212106 367982 0 instr_read_data0\[23\]
rlabel metal2 292622 279956 292622 279956 0 instr_read_data0\[24\]
rlabel metal2 295566 279956 295566 279956 0 instr_read_data0\[25\]
rlabel metal3 133653 476204 133653 476204 0 instr_read_data0\[26\]
rlabel metal3 136229 476204 136229 476204 0 instr_read_data0\[27\]
rlabel metal3 138897 476204 138897 476204 0 instr_read_data0\[28\]
rlabel metal3 141565 476204 141565 476204 0 instr_read_data0\[29\]
rlabel metal2 217826 279956 217826 279956 0 instr_read_data0\[2\]
rlabel metal2 310286 279956 310286 279956 0 instr_read_data0\[30\]
rlabel metal2 313230 279956 313230 279956 0 instr_read_data0\[31\]
rlabel metal3 76659 476204 76659 476204 0 instr_read_data0\[3\]
rlabel metal3 78545 476204 78545 476204 0 instr_read_data0\[4\]
rlabel metal2 230706 279956 230706 279956 0 instr_read_data0\[5\]
rlabel metal2 234846 279956 234846 279956 0 instr_read_data0\[6\]
rlabel metal1 146832 448018 146832 448018 0 instr_read_data0\[7\]
rlabel metal1 147476 448086 147476 448086 0 instr_read_data0\[8\]
rlabel metal1 148810 448154 148810 448154 0 instr_read_data0\[9\]
rlabel metal3 68655 597516 68655 597516 0 instr_read_data1\[0\]
rlabel metal2 249566 279956 249566 279956 0 instr_read_data1\[10\]
rlabel metal2 96554 596343 96554 596343 0 instr_read_data1\[11\]
rlabel metal2 99314 596377 99314 596377 0 instr_read_data1\[12\]
rlabel metal2 102074 596547 102074 596547 0 instr_read_data1\[13\]
rlabel metal4 103316 598128 103316 598128 0 instr_read_data1\[14\]
rlabel metal2 177790 445026 177790 445026 0 instr_read_data1\[15\]
rlabel metal2 180090 444244 180090 444244 0 instr_read_data1\[16\]
rlabel metal2 177882 445876 177882 445876 0 instr_read_data1\[17\]
rlabel metal2 114494 596989 114494 596989 0 instr_read_data1\[18\]
rlabel metal2 117254 597091 117254 597091 0 instr_read_data1\[19\]
rlabel metal2 213778 279956 213778 279956 0 instr_read_data1\[1\]
rlabel via2 118634 596955 118634 596955 0 instr_read_data1\[20\]
rlabel metal2 121394 597125 121394 597125 0 instr_read_data1\[21\]
rlabel metal4 122636 598468 122636 598468 0 instr_read_data1\[22\]
rlabel metal2 177974 446624 177974 446624 0 instr_read_data1\[23\]
rlabel metal2 292990 279956 292990 279956 0 instr_read_data1\[24\]
rlabel metal2 295934 279956 295934 279956 0 instr_read_data1\[25\]
rlabel metal3 133653 597516 133653 597516 0 instr_read_data1\[26\]
rlabel metal3 136229 597516 136229 597516 0 instr_read_data1\[27\]
rlabel via2 139334 597091 139334 597091 0 instr_read_data1\[28\]
rlabel metal3 141565 597516 141565 597516 0 instr_read_data1\[29\]
rlabel metal2 218392 279956 218392 279956 0 instr_read_data1\[2\]
rlabel metal4 141956 598196 141956 598196 0 instr_read_data1\[30\]
rlabel metal2 313598 279956 313598 279956 0 instr_read_data1\[31\]
rlabel metal3 76659 597516 76659 597516 0 instr_read_data1\[3\]
rlabel metal3 78545 597516 78545 597516 0 instr_read_data1\[4\]
rlabel metal3 81213 597516 81213 597516 0 instr_read_data1\[5\]
rlabel metal3 83881 596428 83881 596428 0 instr_read_data1\[6\]
rlabel metal3 86457 597516 86457 597516 0 instr_read_data1\[7\]
rlabel via3 88251 597516 88251 597516 0 instr_read_data1\[8\]
rlabel metal2 91034 596241 91034 596241 0 instr_read_data1\[9\]
rlabel metal2 209822 279956 209822 279956 0 instr_read_data2\[0\]
rlabel metal2 249934 279956 249934 279956 0 instr_read_data2\[10\]
rlabel metal2 253246 279956 253246 279956 0 instr_read_data2\[11\]
rlabel metal2 256558 279956 256558 279956 0 instr_read_data2\[12\]
rlabel metal1 270020 315350 270020 315350 0 instr_read_data2\[13\]
rlabel metal2 263182 279956 263182 279956 0 instr_read_data2\[14\]
rlabel metal1 276092 292026 276092 292026 0 instr_read_data2\[15\]
rlabel metal2 269806 279956 269806 279956 0 instr_read_data2\[16\]
rlabel metal2 272750 279956 272750 279956 0 instr_read_data2\[17\]
rlabel metal2 275694 279956 275694 279956 0 instr_read_data2\[18\]
rlabel metal3 295665 357340 295665 357340 0 instr_read_data2\[19\]
rlabel metal2 214238 279956 214238 279956 0 instr_read_data2\[1\]
rlabel metal1 289892 296106 289892 296106 0 instr_read_data2\[20\]
rlabel metal1 292698 329154 292698 329154 0 instr_read_data2\[21\]
rlabel metal2 287470 279956 287470 279956 0 instr_read_data2\[22\]
rlabel metal2 290414 279956 290414 279956 0 instr_read_data2\[23\]
rlabel metal2 293358 279956 293358 279956 0 instr_read_data2\[24\]
rlabel metal2 296302 279956 296302 279956 0 instr_read_data2\[25\]
rlabel metal3 313375 357340 313375 357340 0 instr_read_data2\[26\]
rlabel metal3 315215 357340 315215 357340 0 instr_read_data2\[27\]
rlabel metal2 305134 279956 305134 279956 0 instr_read_data2\[28\]
rlabel metal2 308078 279956 308078 279956 0 instr_read_data2\[29\]
rlabel metal2 218654 279956 218654 279956 0 instr_read_data2\[2\]
rlabel metal2 311022 279956 311022 279956 0 instr_read_data2\[30\]
rlabel metal2 313966 279956 313966 279956 0 instr_read_data2\[31\]
rlabel metal3 255737 357340 255737 357340 0 instr_read_data2\[3\]
rlabel metal2 227486 279956 227486 279956 0 instr_read_data2\[4\]
rlabel metal2 231534 279956 231534 279956 0 instr_read_data2\[5\]
rlabel metal2 235582 279956 235582 279956 0 instr_read_data2\[6\]
rlabel metal2 239630 279956 239630 279956 0 instr_read_data2\[7\]
rlabel metal3 268065 357340 268065 357340 0 instr_read_data2\[8\]
rlabel metal3 270779 357340 270779 357340 0 instr_read_data2\[9\]
rlabel metal2 210190 279956 210190 279956 0 instr_read_data3\[0\]
rlabel metal2 250302 279956 250302 279956 0 instr_read_data3\[10\]
rlabel metal2 253614 279956 253614 279956 0 instr_read_data3\[11\]
rlabel metal2 214866 416806 214866 416806 0 instr_read_data3\[12\]
rlabel metal2 213118 416874 213118 416874 0 instr_read_data3\[13\]
rlabel metal2 263550 279956 263550 279956 0 instr_read_data3\[14\]
rlabel metal2 266862 279956 266862 279956 0 instr_read_data3\[15\]
rlabel metal2 270174 279956 270174 279956 0 instr_read_data3\[16\]
rlabel metal2 210358 416840 210358 416840 0 instr_read_data3\[17\]
rlabel metal2 276062 279956 276062 279956 0 instr_read_data3\[18\]
rlabel metal2 296286 476153 296286 476153 0 instr_read_data3\[19\]
rlabel metal2 214606 279956 214606 279956 0 instr_read_data3\[1\]
rlabel metal2 281950 279956 281950 279956 0 instr_read_data3\[20\]
rlabel metal2 284894 279956 284894 279956 0 instr_read_data3\[21\]
rlabel metal2 287838 279956 287838 279956 0 instr_read_data3\[22\]
rlabel metal2 290782 279956 290782 279956 0 instr_read_data3\[23\]
rlabel metal2 293726 279956 293726 279956 0 instr_read_data3\[24\]
rlabel metal2 296654 319107 296654 319107 0 instr_read_data3\[25\]
rlabel via2 314594 476595 314594 476595 0 instr_read_data3\[26\]
rlabel metal2 315974 476697 315974 476697 0 instr_read_data3\[27\]
rlabel metal2 305502 279956 305502 279956 0 instr_read_data3\[28\]
rlabel metal2 308446 279956 308446 279956 0 instr_read_data3\[29\]
rlabel metal2 219022 279956 219022 279956 0 instr_read_data3\[2\]
rlabel metal2 311390 279956 311390 279956 0 instr_read_data3\[30\]
rlabel metal2 314334 279956 314334 279956 0 instr_read_data3\[31\]
rlabel metal2 255346 475524 255346 475524 0 instr_read_data3\[3\]
rlabel metal2 227854 279956 227854 279956 0 instr_read_data3\[4\]
rlabel metal2 231902 279956 231902 279956 0 instr_read_data3\[5\]
rlabel metal2 235950 279956 235950 279956 0 instr_read_data3\[6\]
rlabel metal2 239998 279956 239998 279956 0 instr_read_data3\[7\]
rlabel metal2 268042 475439 268042 475439 0 instr_read_data3\[8\]
rlabel metal2 270526 475711 270526 475711 0 instr_read_data3\[9\]
rlabel metal2 210664 279956 210664 279956 0 instr_read_data4\[0\]
rlabel metal4 273516 598400 273516 598400 0 instr_read_data4\[10\]
rlabel metal2 270434 597244 270434 597244 0 instr_read_data4\[11\]
rlabel metal2 277334 598264 277334 598264 0 instr_read_data4\[12\]
rlabel metal2 212382 476901 212382 476901 0 instr_read_data4\[13\]
rlabel metal3 217971 474708 217971 474708 0 instr_read_data4\[14\]
rlabel metal3 285867 597516 285867 597516 0 instr_read_data4\[15\]
rlabel metal3 287661 597108 287661 597108 0 instr_read_data4\[16\]
rlabel metal3 290421 597516 290421 597516 0 instr_read_data4\[17\]
rlabel metal3 292997 597516 292997 597516 0 instr_read_data4\[18\]
rlabel metal2 296378 596241 296378 596241 0 instr_read_data4\[19\]
rlabel metal3 250263 597516 250263 597516 0 instr_read_data4\[1\]
rlabel metal4 298540 598332 298540 598332 0 instr_read_data4\[20\]
rlabel metal4 300932 598400 300932 598400 0 instr_read_data4\[21\]
rlabel metal2 288206 279956 288206 279956 0 instr_read_data4\[22\]
rlabel metal2 291150 279956 291150 279956 0 instr_read_data4\[23\]
rlabel via2 309074 596411 309074 596411 0 instr_read_data4\[24\]
rlabel metal2 311834 596649 311834 596649 0 instr_read_data4\[25\]
rlabel metal2 314594 596649 314594 596649 0 instr_read_data4\[26\]
rlabel via2 315974 596547 315974 596547 0 instr_read_data4\[27\]
rlabel via2 318734 596683 318734 596683 0 instr_read_data4\[28\]
rlabel metal2 308814 279956 308814 279956 0 instr_read_data4\[29\]
rlabel metal4 253644 597924 253644 597924 0 instr_read_data4\[2\]
rlabel metal2 311758 279956 311758 279956 0 instr_read_data4\[30\]
rlabel metal2 327014 596921 327014 596921 0 instr_read_data4\[31\]
rlabel metal4 256036 597992 256036 597992 0 instr_read_data4\[3\]
rlabel metal4 257876 597810 257876 597810 0 instr_read_data4\[4\]
rlabel metal2 213578 477836 213578 477836 0 instr_read_data4\[5\]
rlabel metal2 213670 475184 213670 475184 0 instr_read_data4\[6\]
rlabel metal2 213762 475048 213762 475048 0 instr_read_data4\[7\]
rlabel metal3 268065 597516 268065 597516 0 instr_read_data4\[8\]
rlabel metal3 270733 597516 270733 597516 0 instr_read_data4\[9\]
rlabel metal2 210926 279956 210926 279956 0 instr_read_data5\[0\]
rlabel metal2 251038 279956 251038 279956 0 instr_read_data5\[10\]
rlabel metal2 254350 279956 254350 279956 0 instr_read_data5\[11\]
rlabel metal2 257662 279956 257662 279956 0 instr_read_data5\[12\]
rlabel via2 460966 356099 460966 356099 0 instr_read_data5\[13\]
rlabel metal3 462967 357340 462967 357340 0 instr_read_data5\[14\]
rlabel metal3 465175 357340 465175 357340 0 instr_read_data5\[15\]
rlabel metal2 270910 279956 270910 279956 0 instr_read_data5\[16\]
rlabel metal2 273854 279956 273854 279956 0 instr_read_data5\[17\]
rlabel metal2 276798 279956 276798 279956 0 instr_read_data5\[18\]
rlabel metal2 467222 332350 467222 332350 0 instr_read_data5\[19\]
rlabel metal2 215342 279956 215342 279956 0 instr_read_data5\[1\]
rlabel metal1 376970 307054 376970 307054 0 instr_read_data5\[20\]
rlabel metal2 480562 356609 480562 356609 0 instr_read_data5\[21\]
rlabel metal2 288574 279956 288574 279956 0 instr_read_data5\[22\]
rlabel metal2 291518 279956 291518 279956 0 instr_read_data5\[23\]
rlabel metal2 294462 279956 294462 279956 0 instr_read_data5\[24\]
rlabel metal4 489716 357816 489716 357816 0 instr_read_data5\[25\]
rlabel metal1 388608 311134 388608 311134 0 instr_read_data5\[26\]
rlabel metal2 487830 332962 487830 332962 0 instr_read_data5\[27\]
rlabel metal2 306238 279956 306238 279956 0 instr_read_data5\[28\]
rlabel metal2 309182 279956 309182 279956 0 instr_read_data5\[29\]
rlabel metal2 219758 279956 219758 279956 0 instr_read_data5\[2\]
rlabel metal2 312126 279956 312126 279956 0 instr_read_data5\[30\]
rlabel metal2 315070 279956 315070 279956 0 instr_read_data5\[31\]
rlabel metal1 329452 331874 329452 331874 0 instr_read_data5\[3\]
rlabel metal2 228590 279956 228590 279956 0 instr_read_data5\[4\]
rlabel metal2 232638 279956 232638 279956 0 instr_read_data5\[5\]
rlabel metal2 236686 279956 236686 279956 0 instr_read_data5\[6\]
rlabel via3 445901 357340 445901 357340 0 instr_read_data5\[7\]
rlabel metal3 447787 357340 447787 357340 0 instr_read_data5\[8\]
rlabel metal3 450501 357340 450501 357340 0 instr_read_data5\[9\]
rlabel metal2 211446 279956 211446 279956 0 instr_read_data6\[0\]
rlabel metal2 251406 279956 251406 279956 0 instr_read_data6\[10\]
rlabel metal2 254718 279956 254718 279956 0 instr_read_data6\[11\]
rlabel metal2 258014 317084 258014 317084 0 instr_read_data6\[12\]
rlabel metal4 461012 478516 461012 478516 0 instr_read_data6\[13\]
rlabel metal2 462346 475796 462346 475796 0 instr_read_data6\[14\]
rlabel metal2 267966 279956 267966 279956 0 instr_read_data6\[15\]
rlabel metal2 271278 279956 271278 279956 0 instr_read_data6\[16\]
rlabel metal2 274222 279956 274222 279956 0 instr_read_data6\[17\]
rlabel metal2 277166 279956 277166 279956 0 instr_read_data6\[18\]
rlabel metal2 280110 279956 280110 279956 0 instr_read_data6\[19\]
rlabel metal2 215816 279956 215816 279956 0 instr_read_data6\[1\]
rlabel metal1 339250 354042 339250 354042 0 instr_read_data6\[20\]
rlabel metal2 480562 475405 480562 475405 0 instr_read_data6\[21\]
rlabel metal2 288942 279956 288942 279956 0 instr_read_data6\[22\]
rlabel metal2 291886 279956 291886 279956 0 instr_read_data6\[23\]
rlabel metal2 294830 279956 294830 279956 0 instr_read_data6\[24\]
rlabel metal1 346840 354382 346840 354382 0 instr_read_data6\[25\]
rlabel metal2 300718 279956 300718 279956 0 instr_read_data6\[26\]
rlabel metal2 392426 414290 392426 414290 0 instr_read_data6\[27\]
rlabel metal2 306606 279956 306606 279956 0 instr_read_data6\[28\]
rlabel metal2 309550 279956 309550 279956 0 instr_read_data6\[29\]
rlabel metal3 309465 311100 309465 311100 0 instr_read_data6\[2\]
rlabel metal2 312494 279956 312494 279956 0 instr_read_data6\[30\]
rlabel metal2 315438 279956 315438 279956 0 instr_read_data6\[31\]
rlabel metal2 370530 394859 370530 394859 0 instr_read_data6\[3\]
rlabel metal2 228958 279956 228958 279956 0 instr_read_data6\[4\]
rlabel metal2 233006 279956 233006 279956 0 instr_read_data6\[5\]
rlabel metal2 237054 279956 237054 279956 0 instr_read_data6\[6\]
rlabel metal2 392518 411332 392518 411332 0 instr_read_data6\[7\]
rlabel metal2 393254 411332 393254 411332 0 instr_read_data6\[8\]
rlabel metal2 392794 411332 392794 411332 0 instr_read_data6\[9\]
rlabel metal3 428053 596700 428053 596700 0 instr_read_data7\[0\]
rlabel metal3 446414 596496 446414 596496 0 instr_read_data7\[10\]
rlabel metal2 255086 279956 255086 279956 0 instr_read_data7\[11\]
rlabel metal4 458436 598196 458436 598196 0 instr_read_data7\[12\]
rlabel metal4 461012 598332 461012 598332 0 instr_read_data7\[13\]
rlabel metal3 462967 597516 462967 597516 0 instr_read_data7\[14\]
rlabel metal3 465543 597516 465543 597516 0 instr_read_data7\[15\]
rlabel metal3 468027 597516 468027 597516 0 instr_read_data7\[16\]
rlabel metal4 470396 597856 470396 597856 0 instr_read_data7\[17\]
rlabel metal2 390034 472872 390034 472872 0 instr_read_data7\[18\]
rlabel metal2 390402 472940 390402 472940 0 instr_read_data7\[19\]
rlabel via3 430629 597516 430629 597516 0 instr_read_data7\[1\]
rlabel metal2 390218 472940 390218 472940 0 instr_read_data7\[20\]
rlabel metal3 480585 596972 480585 596972 0 instr_read_data7\[21\]
rlabel metal3 483253 597516 483253 597516 0 instr_read_data7\[22\]
rlabel metal3 485921 597516 485921 597516 0 instr_read_data7\[23\]
rlabel via3 488589 597516 488589 597516 0 instr_read_data7\[24\]
rlabel metal4 489716 597856 489716 597856 0 instr_read_data7\[25\]
rlabel metal2 387458 471682 387458 471682 0 instr_read_data7\[26\]
rlabel metal2 387274 471682 387274 471682 0 instr_read_data7\[27\]
rlabel metal2 306974 279956 306974 279956 0 instr_read_data7\[28\]
rlabel via3 500963 597516 500963 597516 0 instr_read_data7\[29\]
rlabel metal3 326577 563652 326577 563652 0 instr_read_data7\[2\]
rlabel metal3 502849 596972 502849 596972 0 instr_read_data7\[30\]
rlabel metal3 505517 596836 505517 596836 0 instr_read_data7\[31\]
rlabel metal2 434746 597397 434746 597397 0 instr_read_data7\[3\]
rlabel metal2 229326 279956 229326 279956 0 instr_read_data7\[4\]
rlabel metal2 233374 279956 233374 279956 0 instr_read_data7\[5\]
rlabel metal3 443279 597516 443279 597516 0 instr_read_data7\[6\]
rlabel metal3 445855 597516 445855 597516 0 instr_read_data7\[7\]
rlabel metal3 447741 597516 447741 597516 0 instr_read_data7\[8\]
rlabel metal3 450501 597516 450501 597516 0 instr_read_data7\[9\]
rlabel metal2 39790 485180 39790 485180 0 instr_wmask\[0\]
rlabel metal1 39376 485282 39376 485282 0 instr_wmask\[1\]
rlabel metal4 60628 598332 60628 598332 0 instr_wmask\[2\]
rlabel metal2 56442 597312 56442 597312 0 instr_wmask\[3\]
rlabel metal4 63158 599745 63158 599745 0 instr_write_data\[0\]
rlabel metal2 74934 597312 74934 597312 0 instr_write_data\[10\]
rlabel metal4 75942 599745 75942 599745 0 instr_write_data\[11\]
rlabel metal2 77142 596734 77142 596734 0 instr_write_data\[12\]
rlabel metal4 78118 599745 78118 599745 0 instr_write_data\[13\]
rlabel metal4 79478 599745 79478 599745 0 instr_write_data\[14\]
rlabel metal3 79764 596904 79764 596904 0 instr_write_data\[15\]
rlabel metal1 39790 485180 39790 485180 0 instr_write_data\[1\]
rlabel metal4 64676 598468 64676 598468 0 instr_write_data\[2\]
rlabel metal4 83996 598128 83996 598128 0 instr_write_data\[3\]
rlabel metal4 427646 599745 427646 599745 0 instr_write_data\[4\]
rlabel metal4 248734 599813 248734 599813 0 instr_write_data\[5\]
rlabel metal4 250094 599813 250094 599813 0 instr_write_data\[6\]
rlabel metal3 251827 596836 251827 596836 0 instr_write_data\[7\]
rlabel metal4 252406 599813 252406 599813 0 instr_write_data\[8\]
rlabel metal1 249964 350506 249964 350506 0 instr_write_data\[9\]
rlabel metal3 40020 489938 40020 489938 0 instrw_enb
rlabel metal3 581770 6596 581770 6596 0 io_in[0]
rlabel metal2 134902 279956 134902 279956 0 io_in[10]
rlabel metal2 136006 279956 136006 279956 0 io_in[11]
rlabel metal2 579922 563703 579922 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel metal2 139166 279956 139166 279956 0 io_in[14]
rlabel metal2 140270 279956 140270 279956 0 io_in[15]
rlabel metal2 141374 279956 141374 279956 0 io_in[16]
rlabel metal2 392610 521016 392610 521016 0 io_in[17]
rlabel metal2 364366 516467 364366 516467 0 io_in[18]
rlabel metal3 258037 700468 258037 700468 0 io_in[19]
rlabel metal2 121302 164254 121302 164254 0 io_in[1]
rlabel metal4 214452 514216 214452 514216 0 io_in[20]
rlabel metal2 178342 529448 178342 529448 0 io_in[21]
rlabel metal2 178250 491436 178250 491436 0 io_in[22]
rlabel metal2 40020 443292 40020 443292 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 1556 632060 1556 632060 0 io_in[25]
rlabel metal3 1556 579972 1556 579972 0 io_in[26]
rlabel metal3 1878 527884 1878 527884 0 io_in[27]
rlabel metal3 1694 475660 1694 475660 0 io_in[28]
rlabel metal3 1924 423572 1924 423572 0 io_in[29]
rlabel metal2 538982 185130 538982 185130 0 io_in[2]
rlabel metal3 1832 371348 1832 371348 0 io_in[30]
rlabel metal3 1832 319260 1832 319260 0 io_in[31]
rlabel metal3 1832 267172 1832 267172 0 io_in[32]
rlabel metal3 1694 214948 1694 214948 0 io_in[33]
rlabel metal3 1694 162860 1694 162860 0 io_in[34]
rlabel metal3 1832 110636 1832 110636 0 io_in[35]
rlabel metal3 1970 71604 1970 71604 0 io_in[36]
rlabel metal3 1878 32436 1878 32436 0 io_in[37]
rlabel metal2 540270 205088 540270 205088 0 io_in[3]
rlabel metal2 543122 225046 543122 225046 0 io_in[4]
rlabel metal2 544410 245004 544410 245004 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 580198 298435 580198 298435 0 io_in[7]
rlabel via2 580198 351917 580198 351917 0 io_in[8]
rlabel metal2 580198 404651 580198 404651 0 io_in[9]
rlabel metal3 583556 32368 583556 32368 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 136374 279956 136374 279956 0 io_oeb[11]
rlabel metal2 137326 279956 137326 279956 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 140638 279956 140638 279956 0 io_oeb[15]
rlabel metal2 141742 279956 141742 279956 0 io_oeb[16]
rlabel via3 397509 699788 397509 699788 0 io_oeb[17]
rlabel metal4 213164 518840 213164 518840 0 io_oeb[18]
rlabel metal4 211692 521764 211692 521764 0 io_oeb[19]
rlabel metal2 538982 78657 538982 78657 0 io_oeb[1]
rlabel metal2 146158 279820 146158 279820 0 io_oeb[20]
rlabel metal2 137862 702076 137862 702076 0 io_oeb[21]
rlabel metal2 178158 491589 178158 491589 0 io_oeb[22]
rlabel metal1 78200 313922 78200 313922 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 1786 606084 1786 606084 0 io_oeb[25]
rlabel metal3 1878 553860 1878 553860 0 io_oeb[26]
rlabel metal3 1694 501772 1694 501772 0 io_oeb[27]
rlabel metal3 1740 449548 1740 449548 0 io_oeb[28]
rlabel metal3 1832 397460 1832 397460 0 io_oeb[29]
rlabel metal2 543030 198050 543030 198050 0 io_oeb[2]
rlabel metal3 1832 345372 1832 345372 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 1832 241060 1832 241060 0 io_oeb[32]
rlabel metal3 1832 188836 1832 188836 0 io_oeb[33]
rlabel metal3 1832 136748 1832 136748 0 io_oeb[34]
rlabel metal3 2016 84660 2016 84660 0 io_oeb[35]
rlabel metal3 1924 45492 1924 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal3 581954 152660 581954 152660 0 io_oeb[3]
rlabel metal3 582092 192508 582092 192508 0 io_oeb[4]
rlabel metal2 580014 232781 580014 232781 0 io_oeb[5]
rlabel metal3 442727 271932 442727 271932 0 io_oeb[6]
rlabel metal2 580198 324785 580198 324785 0 io_oeb[7]
rlabel metal2 132910 279956 132910 279956 0 io_oeb[8]
rlabel metal2 580198 431103 580198 431103 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 135486 279956 135486 279956 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal2 579646 577269 579646 577269 0 io_out[12]
rlabel metal2 138798 279956 138798 279956 0 io_out[13]
rlabel metal2 139902 279956 139902 279956 0 io_out[14]
rlabel metal2 141006 279956 141006 279956 0 io_out[15]
rlabel metal2 142094 299693 142094 299693 0 io_out[16]
rlabel metal2 366390 512686 366390 512686 0 io_out[17]
rlabel metal2 177330 492762 177330 492762 0 io_out[18]
rlabel metal2 177422 492864 177422 492864 0 io_out[19]
rlabel metal3 581908 59636 581908 59636 0 io_out[1]
rlabel metal2 219006 701974 219006 701974 0 io_out[20]
rlabel metal2 154146 702110 154146 702110 0 io_out[21]
rlabel metal2 176686 491368 176686 491368 0 io_out[22]
rlabel metal2 24334 701634 24334 701634 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal2 3496 306360 3496 306360 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 1924 410516 1924 410516 0 io_out[29]
rlabel metal3 582000 99484 582000 99484 0 io_out[2]
rlabel metal3 1832 358428 1832 358428 0 io_out[30]
rlabel metal3 1878 306204 1878 306204 0 io_out[31]
rlabel metal3 1648 254116 1648 254116 0 io_out[32]
rlabel metal3 2062 201892 2062 201892 0 io_out[33]
rlabel metal3 1832 149804 1832 149804 0 io_out[34]
rlabel metal3 1832 97580 1832 97580 0 io_out[35]
rlabel metal3 1924 58548 1924 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 579830 139349 579830 139349 0 io_out[3]
rlabel metal3 582046 179180 582046 179180 0 io_out[4]
rlabel metal3 582138 219028 582138 219028 0 io_out[5]
rlabel metal2 579830 259131 579830 259131 0 io_out[6]
rlabel metal2 580198 311967 580198 311967 0 io_out[7]
rlabel metal2 579830 364735 579830 364735 0 io_out[8]
rlabel metal2 134382 279956 134382 279956 0 io_out[9]
rlabel metal2 125757 340 125757 340 0 la_data_in[0]
rlabel metal2 127298 80036 127298 80036 0 la_data_out[0]
rlabel metal2 481712 16560 481712 16560 0 la_data_out[100]
rlabel metal2 485017 340 485017 340 0 la_data_out[101]
rlabel metal2 268012 80036 268012 80036 0 la_data_out[102]
rlabel metal2 269392 80036 269392 80036 0 la_data_out[103]
rlabel metal2 270772 80036 270772 80036 0 la_data_out[104]
rlabel metal2 272152 80036 272152 80036 0 la_data_out[105]
rlabel metal2 273532 80036 273532 80036 0 la_data_out[106]
rlabel metal2 274912 80036 274912 80036 0 la_data_out[107]
rlabel metal2 276292 80036 276292 80036 0 la_data_out[108]
rlabel metal2 277672 80036 277672 80036 0 la_data_out[109]
rlabel metal2 141052 80036 141052 80036 0 la_data_out[10]
rlabel metal2 279052 80036 279052 80036 0 la_data_out[110]
rlabel metal2 520766 2812 520766 2812 0 la_data_out[111]
rlabel metal2 524262 2778 524262 2778 0 la_data_out[112]
rlabel metal2 527850 2744 527850 2744 0 la_data_out[113]
rlabel metal2 284572 80036 284572 80036 0 la_data_out[114]
rlabel metal2 285952 80036 285952 80036 0 la_data_out[115]
rlabel metal2 287332 80036 287332 80036 0 la_data_out[116]
rlabel metal2 288712 80036 288712 80036 0 la_data_out[117]
rlabel metal2 290092 80036 290092 80036 0 la_data_out[118]
rlabel metal2 291472 80036 291472 80036 0 la_data_out[119]
rlabel metal2 142432 80036 142432 80036 0 la_data_out[11]
rlabel metal2 292852 80036 292852 80036 0 la_data_out[120]
rlabel metal2 294232 80036 294232 80036 0 la_data_out[121]
rlabel metal2 295612 80036 295612 80036 0 la_data_out[122]
rlabel metal2 563171 340 563171 340 0 la_data_out[123]
rlabel metal2 565846 21047 565846 21047 0 la_data_out[124]
rlabel metal2 299752 80036 299752 80036 0 la_data_out[125]
rlabel metal2 301132 80036 301132 80036 0 la_data_out[126]
rlabel metal2 577201 340 577201 340 0 la_data_out[127]
rlabel metal2 143812 80036 143812 80036 0 la_data_out[12]
rlabel metal2 173190 2098 173190 2098 0 la_data_out[13]
rlabel metal2 176686 2064 176686 2064 0 la_data_out[14]
rlabel metal2 180274 2030 180274 2030 0 la_data_out[15]
rlabel metal2 149332 80036 149332 80036 0 la_data_out[16]
rlabel metal2 150712 80036 150712 80036 0 la_data_out[17]
rlabel metal2 152092 80036 152092 80036 0 la_data_out[18]
rlabel metal2 153472 80036 153472 80036 0 la_data_out[19]
rlabel metal2 130594 1911 130594 1911 0 la_data_out[1]
rlabel metal1 156032 77282 156032 77282 0 la_data_out[20]
rlabel metal1 157412 77282 157412 77282 0 la_data_out[21]
rlabel metal1 158792 77282 158792 77282 0 la_data_out[22]
rlabel metal2 159574 79101 159574 79101 0 la_data_out[23]
rlabel metal2 160954 79067 160954 79067 0 la_data_out[24]
rlabel metal2 215503 340 215503 340 0 la_data_out[25]
rlabel metal2 219282 1894 219282 1894 0 la_data_out[26]
rlabel metal2 165094 77605 165094 77605 0 la_data_out[27]
rlabel metal2 165892 80036 165892 80036 0 la_data_out[28]
rlabel metal2 229625 340 229625 340 0 la_data_out[29]
rlabel metal2 134182 2234 134182 2234 0 la_data_out[2]
rlabel metal2 233358 16560 233358 16560 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal1 172592 77282 172592 77282 0 la_data_out[32]
rlabel metal2 172792 80036 172792 80036 0 la_data_out[33]
rlabel metal2 174172 80036 174172 80036 0 la_data_out[34]
rlabel metal2 175552 80036 175552 80036 0 la_data_out[35]
rlabel metal2 176932 80036 176932 80036 0 la_data_out[36]
rlabel metal2 178312 80036 178312 80036 0 la_data_out[37]
rlabel metal2 179692 80036 179692 80036 0 la_data_out[38]
rlabel metal2 181072 80036 181072 80036 0 la_data_out[39]
rlabel metal2 137678 1996 137678 1996 0 la_data_out[3]
rlabel metal2 268870 2676 268870 2676 0 la_data_out[40]
rlabel metal2 272458 2642 272458 2642 0 la_data_out[41]
rlabel metal2 276046 2608 276046 2608 0 la_data_out[42]
rlabel metal2 186592 80036 186592 80036 0 la_data_out[43]
rlabel metal2 199410 41038 199410 41038 0 la_data_out[44]
rlabel metal2 189934 79271 189934 79271 0 la_data_out[45]
rlabel metal2 191314 79237 191314 79237 0 la_data_out[46]
rlabel metal2 192694 79203 192694 79203 0 la_data_out[47]
rlabel metal2 194074 79135 194074 79135 0 la_data_out[48]
rlabel metal2 195454 79169 195454 79169 0 la_data_out[49]
rlabel metal2 141266 1894 141266 1894 0 la_data_out[4]
rlabel metal2 196252 80036 196252 80036 0 la_data_out[50]
rlabel metal2 197632 80036 197632 80036 0 la_data_out[51]
rlabel metal2 199012 80036 199012 80036 0 la_data_out[52]
rlabel metal2 315054 3526 315054 3526 0 la_data_out[53]
rlabel metal2 201772 80036 201772 80036 0 la_data_out[54]
rlabel metal2 203152 80036 203152 80036 0 la_data_out[55]
rlabel metal2 204532 80036 204532 80036 0 la_data_out[56]
rlabel metal2 329222 3390 329222 3390 0 la_data_out[57]
rlabel metal2 332718 3356 332718 3356 0 la_data_out[58]
rlabel metal2 208718 80036 208718 80036 0 la_data_out[59]
rlabel metal2 134198 80036 134198 80036 0 la_data_out[5]
rlabel metal2 210052 80036 210052 80036 0 la_data_out[60]
rlabel metal2 211478 80036 211478 80036 0 la_data_out[61]
rlabel metal2 212812 80036 212812 80036 0 la_data_out[62]
rlabel metal1 216062 77282 216062 77282 0 la_data_out[63]
rlabel metal2 215618 80036 215618 80036 0 la_data_out[64]
rlabel metal2 216952 80036 216952 80036 0 la_data_out[65]
rlabel metal2 218914 78999 218914 78999 0 la_data_out[66]
rlabel metal2 364366 19007 364366 19007 0 la_data_out[67]
rlabel metal2 367993 340 367993 340 0 la_data_out[68]
rlabel metal2 371489 340 371489 340 0 la_data_out[69]
rlabel metal1 138322 3502 138322 3502 0 la_data_out[6]
rlabel metal2 223852 80036 223852 80036 0 la_data_out[70]
rlabel metal2 231150 52802 231150 52802 0 la_data_out[71]
rlabel metal2 226612 80036 226612 80036 0 la_data_out[72]
rlabel metal2 385526 16560 385526 16560 0 la_data_out[73]
rlabel metal2 229372 80036 229372 80036 0 la_data_out[74]
rlabel metal2 230752 80036 230752 80036 0 la_data_out[75]
rlabel metal2 232132 80036 232132 80036 0 la_data_out[76]
rlabel metal2 234094 79339 234094 79339 0 la_data_out[77]
rlabel metal2 234892 80036 234892 80036 0 la_data_out[78]
rlabel metal2 236854 79033 236854 79033 0 la_data_out[79]
rlabel metal2 136912 80036 136912 80036 0 la_data_out[7]
rlabel metal2 237652 80036 237652 80036 0 la_data_out[80]
rlabel metal1 242282 77418 242282 77418 0 la_data_out[81]
rlabel metal1 241638 77282 241638 77282 0 la_data_out[82]
rlabel metal1 244352 77350 244352 77350 0 la_data_out[83]
rlabel metal2 424994 4172 424994 4172 0 la_data_out[84]
rlabel metal2 427846 16933 427846 16933 0 la_data_out[85]
rlabel metal2 245932 80036 245932 80036 0 la_data_out[86]
rlabel metal2 313950 40868 313950 40868 0 la_data_out[87]
rlabel metal2 248692 80036 248692 80036 0 la_data_out[88]
rlabel metal2 250072 80036 250072 80036 0 la_data_out[89]
rlabel metal2 138292 80036 138292 80036 0 la_data_out[8]
rlabel metal2 251452 80036 251452 80036 0 la_data_out[90]
rlabel metal2 252832 80036 252832 80036 0 la_data_out[91]
rlabel metal2 254212 80036 254212 80036 0 la_data_out[92]
rlabel metal2 256174 79033 256174 79033 0 la_data_out[93]
rlabel metal2 256972 80036 256972 80036 0 la_data_out[94]
rlabel metal2 464002 8150 464002 8150 0 la_data_out[95]
rlabel metal2 467498 4002 467498 4002 0 la_data_out[96]
rlabel metal2 261694 79067 261694 79067 0 la_data_out[97]
rlabel metal2 262492 80036 262492 80036 0 la_data_out[98]
rlabel metal2 263872 80036 263872 80036 0 la_data_out[99]
rlabel metal2 139672 80036 139672 80036 0 la_data_out[9]
rlabel metal2 128202 1894 128202 1894 0 la_oenb[0]
rlabel metal1 178802 444346 178802 444346 0 low
rlabel metal2 309412 80036 309412 80036 0 reset
rlabel metal2 311374 79237 311374 79237 0 start
rlabel metal2 178066 281758 178066 281758 0 uP_data_mem_addr\[0\]
rlabel metal2 434187 229908 434187 229908 0 uP_data_mem_addr\[1\]
rlabel metal2 436579 229908 436579 229908 0 uP_data_mem_addr\[2\]
rlabel metal2 171702 279956 171702 279956 0 uP_data_mem_addr\[3\]
rlabel metal2 173542 279956 173542 279956 0 uP_data_mem_addr\[4\]
rlabel metal2 443755 229908 443755 229908 0 uP_data_mem_addr\[5\]
rlabel metal2 446147 229908 446147 229908 0 uP_data_mem_addr\[6\]
rlabel metal2 448631 229908 448631 229908 0 uP_data_mem_addr\[7\]
rlabel metal2 527666 231258 527666 231258 0 uP_dataw_en
rlabel metal2 179446 280670 179446 280670 0 uP_instr\[0\]
rlabel metal2 410267 229908 410267 229908 0 uP_instr\[10\]
rlabel metal2 415051 229908 415051 229908 0 uP_instr\[11\]
rlabel metal2 419835 229908 419835 229908 0 uP_instr\[12\]
rlabel metal2 424619 229908 424619 229908 0 uP_instr\[13\]
rlabel metal2 427011 229908 427011 229908 0 uP_instr\[14\]
rlabel metal2 429403 229908 429403 229908 0 uP_instr\[15\]
rlabel metal2 367257 229908 367257 229908 0 uP_instr\[1\]
rlabel metal2 371995 229908 371995 229908 0 uP_instr\[2\]
rlabel metal2 172070 279956 172070 279956 0 uP_instr\[3\]
rlabel metal2 173758 279956 173758 279956 0 uP_instr\[4\]
rlabel metal2 386485 229908 386485 229908 0 uP_instr\[5\]
rlabel metal2 391131 229908 391131 229908 0 uP_instr\[6\]
rlabel metal2 179278 279820 179278 279820 0 uP_instr\[7\]
rlabel metal2 180734 280245 180734 280245 0 uP_instr\[8\]
rlabel metal2 405483 229908 405483 229908 0 uP_instr\[9\]
rlabel metal2 364819 229908 364819 229908 0 uP_instr_mem_addr\[0\]
rlabel metal2 412751 229908 412751 229908 0 uP_instr_mem_addr\[10\]
rlabel metal2 417443 229908 417443 229908 0 uP_instr_mem_addr\[11\]
rlabel metal2 422365 229908 422365 229908 0 uP_instr_mem_addr\[12\]
rlabel metal2 369603 229908 369603 229908 0 uP_instr_mem_addr\[1\]
rlabel metal2 374387 229908 374387 229908 0 uP_instr_mem_addr\[2\]
rlabel metal2 172392 279956 172392 279956 0 uP_instr_mem_addr\[3\]
rlabel metal2 383955 229908 383955 229908 0 uP_instr_mem_addr\[4\]
rlabel metal2 388739 229908 388739 229908 0 uP_instr_mem_addr\[5\]
rlabel metal2 177912 279956 177912 279956 0 uP_instr_mem_addr\[6\]
rlabel metal2 179798 279956 179798 279956 0 uP_instr_mem_addr\[7\]
rlabel metal2 403137 229908 403137 229908 0 uP_instr_mem_addr\[8\]
rlabel metal2 407875 229908 407875 229908 0 uP_instr_mem_addr\[9\]
rlabel metal2 450931 229908 450931 229908 0 uP_read_data\[0\]
rlabel metal2 474897 229908 474897 229908 0 uP_read_data\[10\]
rlabel metal2 191682 281588 191682 281588 0 uP_read_data\[11\]
rlabel metal2 479635 229908 479635 229908 0 uP_read_data\[12\]
rlabel metal2 482027 229908 482027 229908 0 uP_read_data\[13\]
rlabel metal2 484511 229908 484511 229908 0 uP_read_data\[14\]
rlabel metal2 486811 229908 486811 229908 0 uP_read_data\[15\]
rlabel metal2 453369 229908 453369 229908 0 uP_read_data\[1\]
rlabel metal2 455906 231428 455906 231428 0 uP_read_data\[2\]
rlabel metal2 172654 279956 172654 279956 0 uP_read_data\[3\]
rlabel metal2 174646 279956 174646 279956 0 uP_read_data\[4\]
rlabel metal2 462891 229908 462891 229908 0 uP_read_data\[5\]
rlabel metal2 465474 231938 465474 231938 0 uP_read_data\[6\]
rlabel metal2 180166 279956 180166 279956 0 uP_read_data\[7\]
rlabel metal2 470021 229908 470021 229908 0 uP_read_data\[8\]
rlabel metal2 472459 229908 472459 229908 0 uP_read_data\[9\]
rlabel metal2 489394 231462 489394 231462 0 uP_write_data\[0\]
rlabel metal2 513314 231207 513314 231207 0 uP_write_data\[10\]
rlabel metal2 515515 229908 515515 229908 0 uP_write_data\[11\]
rlabel metal2 517907 229908 517907 229908 0 uP_write_data\[12\]
rlabel metal2 520490 231428 520490 231428 0 uP_write_data\[13\]
rlabel metal2 522882 231224 522882 231224 0 uP_write_data\[14\]
rlabel metal2 525274 231394 525274 231394 0 uP_write_data\[15\]
rlabel metal2 314870 280942 314870 280942 0 uP_write_data\[1\]
rlabel metal2 171334 279956 171334 279956 0 uP_write_data\[2\]
rlabel metal2 173022 279956 173022 279956 0 uP_write_data\[3\]
rlabel metal2 174968 279956 174968 279956 0 uP_write_data\[4\]
rlabel metal2 501354 231326 501354 231326 0 uP_write_data\[5\]
rlabel metal2 503746 231462 503746 231462 0 uP_write_data\[6\]
rlabel metal2 505947 229908 505947 229908 0 uP_write_data\[7\]
rlabel metal2 508530 231292 508530 231292 0 uP_write_data\[8\]
rlabel metal2 510922 231258 510922 231258 0 uP_write_data\[9\]
rlabel metal2 581026 1894 581026 1894 0 user_irq[0]
rlabel metal2 582222 1962 582222 1962 0 user_irq[1]
rlabel metal2 307234 79135 307234 79135 0 user_irq[2]
rlabel metal2 361 340 361 340 0 wb_clk_i
rlabel metal2 1557 340 1557 340 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
