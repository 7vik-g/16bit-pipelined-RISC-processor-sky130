* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for sky130_sram_2kbyte_1rw1r_32x512_8 abstract view
.subckt sky130_sram_2kbyte_1rw1r_32x512_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr1[0]
+ addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] addr1[8] csb0 csb1
+ web0 clk0 clk1 wmask0[0] wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2]
+ dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[30] dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4]
+ dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13]
+ dout1[14] dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[20] dout1[21]
+ dout1[22] dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29]
+ dout1[30] dout1[31] vccd1 vssd1
.ends

* Black-box entry subcircuit for io_interface abstract view
.subckt io_interface Serial_input Serial_output clk data_mem_addr[0] data_mem_addr[1]
+ data_mem_addr[2] data_mem_addr[3] data_mem_addr[4] data_mem_addr[5] data_mem_addr[6]
+ data_mem_addr[7] data_mem_csb data_read_data[0] data_read_data[10] data_read_data[11]
+ data_read_data[12] data_read_data[13] data_read_data[14] data_read_data[15] data_read_data[1]
+ data_read_data[2] data_read_data[3] data_read_data[4] data_read_data[5] data_read_data[6]
+ data_read_data[7] data_read_data[8] data_read_data[9] data_wmask[0] data_wmask[1]
+ data_wmask[2] data_wmask[3] data_write_data[0] data_write_data[10] data_write_data[11]
+ data_write_data[12] data_write_data[13] data_write_data[14] data_write_data[15]
+ data_write_data[1] data_write_data[2] data_write_data[3] data_write_data[4] data_write_data[5]
+ data_write_data[6] data_write_data[7] data_write_data[8] data_write_data[9] dataw_enb
+ high hlt instr_mem_addr_9bit[0] instr_mem_addr_9bit[1] instr_mem_addr_9bit[2] instr_mem_addr_9bit[3]
+ instr_mem_addr_9bit[4] instr_mem_addr_9bit[5] instr_mem_addr_9bit[6] instr_mem_addr_9bit[7]
+ instr_mem_addr_9bit[8] instr_mem_csb[0] instr_mem_csb[1] instr_mem_csb[2] instr_mem_csb[3]
+ instr_mem_csb[4] instr_mem_csb[5] instr_mem_csb[6] instr_mem_csb[7] instr_read_data0[0]
+ instr_read_data0[10] instr_read_data0[11] instr_read_data0[12] instr_read_data0[13]
+ instr_read_data0[14] instr_read_data0[15] instr_read_data0[16] instr_read_data0[17]
+ instr_read_data0[18] instr_read_data0[19] instr_read_data0[1] instr_read_data0[20]
+ instr_read_data0[21] instr_read_data0[22] instr_read_data0[23] instr_read_data0[24]
+ instr_read_data0[25] instr_read_data0[26] instr_read_data0[27] instr_read_data0[28]
+ instr_read_data0[29] instr_read_data0[2] instr_read_data0[30] instr_read_data0[31]
+ instr_read_data0[3] instr_read_data0[4] instr_read_data0[5] instr_read_data0[6]
+ instr_read_data0[7] instr_read_data0[8] instr_read_data0[9] instr_read_data1[0]
+ instr_read_data1[10] instr_read_data1[11] instr_read_data1[12] instr_read_data1[13]
+ instr_read_data1[14] instr_read_data1[15] instr_read_data1[16] instr_read_data1[17]
+ instr_read_data1[18] instr_read_data1[19] instr_read_data1[1] instr_read_data1[20]
+ instr_read_data1[21] instr_read_data1[22] instr_read_data1[23] instr_read_data1[24]
+ instr_read_data1[25] instr_read_data1[26] instr_read_data1[27] instr_read_data1[28]
+ instr_read_data1[29] instr_read_data1[2] instr_read_data1[30] instr_read_data1[31]
+ instr_read_data1[3] instr_read_data1[4] instr_read_data1[5] instr_read_data1[6]
+ instr_read_data1[7] instr_read_data1[8] instr_read_data1[9] instr_read_data2[0]
+ instr_read_data2[10] instr_read_data2[11] instr_read_data2[12] instr_read_data2[13]
+ instr_read_data2[14] instr_read_data2[15] instr_read_data2[16] instr_read_data2[17]
+ instr_read_data2[18] instr_read_data2[19] instr_read_data2[1] instr_read_data2[20]
+ instr_read_data2[21] instr_read_data2[22] instr_read_data2[23] instr_read_data2[24]
+ instr_read_data2[25] instr_read_data2[26] instr_read_data2[27] instr_read_data2[28]
+ instr_read_data2[29] instr_read_data2[2] instr_read_data2[30] instr_read_data2[31]
+ instr_read_data2[3] instr_read_data2[4] instr_read_data2[5] instr_read_data2[6]
+ instr_read_data2[7] instr_read_data2[8] instr_read_data2[9] instr_read_data3[0]
+ instr_read_data3[10] instr_read_data3[11] instr_read_data3[12] instr_read_data3[13]
+ instr_read_data3[14] instr_read_data3[15] instr_read_data3[16] instr_read_data3[17]
+ instr_read_data3[18] instr_read_data3[19] instr_read_data3[1] instr_read_data3[20]
+ instr_read_data3[21] instr_read_data3[22] instr_read_data3[23] instr_read_data3[24]
+ instr_read_data3[25] instr_read_data3[26] instr_read_data3[27] instr_read_data3[28]
+ instr_read_data3[29] instr_read_data3[2] instr_read_data3[30] instr_read_data3[31]
+ instr_read_data3[3] instr_read_data3[4] instr_read_data3[5] instr_read_data3[6]
+ instr_read_data3[7] instr_read_data3[8] instr_read_data3[9] instr_read_data4[0]
+ instr_read_data4[10] instr_read_data4[11] instr_read_data4[12] instr_read_data4[13]
+ instr_read_data4[14] instr_read_data4[15] instr_read_data4[16] instr_read_data4[17]
+ instr_read_data4[18] instr_read_data4[19] instr_read_data4[1] instr_read_data4[20]
+ instr_read_data4[21] instr_read_data4[22] instr_read_data4[23] instr_read_data4[24]
+ instr_read_data4[25] instr_read_data4[26] instr_read_data4[27] instr_read_data4[28]
+ instr_read_data4[29] instr_read_data4[2] instr_read_data4[30] instr_read_data4[31]
+ instr_read_data4[3] instr_read_data4[4] instr_read_data4[5] instr_read_data4[6]
+ instr_read_data4[7] instr_read_data4[8] instr_read_data4[9] instr_read_data5[0]
+ instr_read_data5[10] instr_read_data5[11] instr_read_data5[12] instr_read_data5[13]
+ instr_read_data5[14] instr_read_data5[15] instr_read_data5[16] instr_read_data5[17]
+ instr_read_data5[18] instr_read_data5[19] instr_read_data5[1] instr_read_data5[20]
+ instr_read_data5[21] instr_read_data5[22] instr_read_data5[23] instr_read_data5[24]
+ instr_read_data5[25] instr_read_data5[26] instr_read_data5[27] instr_read_data5[28]
+ instr_read_data5[29] instr_read_data5[2] instr_read_data5[30] instr_read_data5[31]
+ instr_read_data5[3] instr_read_data5[4] instr_read_data5[5] instr_read_data5[6]
+ instr_read_data5[7] instr_read_data5[8] instr_read_data5[9] instr_read_data6[0]
+ instr_read_data6[10] instr_read_data6[11] instr_read_data6[12] instr_read_data6[13]
+ instr_read_data6[14] instr_read_data6[15] instr_read_data6[16] instr_read_data6[17]
+ instr_read_data6[18] instr_read_data6[19] instr_read_data6[1] instr_read_data6[20]
+ instr_read_data6[21] instr_read_data6[22] instr_read_data6[23] instr_read_data6[24]
+ instr_read_data6[25] instr_read_data6[26] instr_read_data6[27] instr_read_data6[28]
+ instr_read_data6[29] instr_read_data6[2] instr_read_data6[30] instr_read_data6[31]
+ instr_read_data6[3] instr_read_data6[4] instr_read_data6[5] instr_read_data6[6]
+ instr_read_data6[7] instr_read_data6[8] instr_read_data6[9] instr_read_data7[0]
+ instr_read_data7[10] instr_read_data7[11] instr_read_data7[12] instr_read_data7[13]
+ instr_read_data7[14] instr_read_data7[15] instr_read_data7[16] instr_read_data7[17]
+ instr_read_data7[18] instr_read_data7[19] instr_read_data7[1] instr_read_data7[20]
+ instr_read_data7[21] instr_read_data7[22] instr_read_data7[23] instr_read_data7[24]
+ instr_read_data7[25] instr_read_data7[26] instr_read_data7[27] instr_read_data7[28]
+ instr_read_data7[29] instr_read_data7[2] instr_read_data7[30] instr_read_data7[31]
+ instr_read_data7[3] instr_read_data7[4] instr_read_data7[5] instr_read_data7[6]
+ instr_read_data7[7] instr_read_data7[8] instr_read_data7[9] instr_wmask[0] instr_wmask[1]
+ instr_wmask[2] instr_wmask[3] instr_write_data[0] instr_write_data[10] instr_write_data[11]
+ instr_write_data[12] instr_write_data[13] instr_write_data[14] instr_write_data[15]
+ instr_write_data[1] instr_write_data[2] instr_write_data[3] instr_write_data[4]
+ instr_write_data[5] instr_write_data[6] instr_write_data[7] instr_write_data[8]
+ instr_write_data[9] instrw_enb io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] irq[0] irq[1] irq[2] la_data_in la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb low reset start uP_data_mem_addr[0]
+ uP_data_mem_addr[1] uP_data_mem_addr[2] uP_data_mem_addr[3] uP_data_mem_addr[4]
+ uP_data_mem_addr[5] uP_data_mem_addr[6] uP_data_mem_addr[7] uP_dataw_en uP_instr[0]
+ uP_instr[10] uP_instr[11] uP_instr[12] uP_instr[13] uP_instr[14] uP_instr[15] uP_instr[1]
+ uP_instr[2] uP_instr[3] uP_instr[4] uP_instr[5] uP_instr[6] uP_instr[7] uP_instr[8]
+ uP_instr[9] uP_instr_mem_addr[0] uP_instr_mem_addr[10] uP_instr_mem_addr[11] uP_instr_mem_addr[12]
+ uP_instr_mem_addr[1] uP_instr_mem_addr[2] uP_instr_mem_addr[3] uP_instr_mem_addr[4]
+ uP_instr_mem_addr[5] uP_instr_mem_addr[6] uP_instr_mem_addr[7] uP_instr_mem_addr[8]
+ uP_instr_mem_addr[9] uP_read_data[0] uP_read_data[10] uP_read_data[11] uP_read_data[12]
+ uP_read_data[13] uP_read_data[14] uP_read_data[15] uP_read_data[1] uP_read_data[2]
+ uP_read_data[3] uP_read_data[4] uP_read_data[5] uP_read_data[6] uP_read_data[7]
+ uP_read_data[8] uP_read_data[9] uP_write_data[0] uP_write_data[10] uP_write_data[11]
+ uP_write_data[12] uP_write_data[13] uP_write_data[14] uP_write_data[15] uP_write_data[1]
+ uP_write_data[2] uP_write_data[3] uP_write_data[4] uP_write_data[5] uP_write_data[6]
+ uP_write_data[7] uP_write_data[8] uP_write_data[9] vccd1 vssd1 wb_clk_i wb_rst_i
.ends

* Black-box entry subcircuit for processor abstract view
.subckt processor Dataw_en Serial_input Serial_output clk data_mem_addr[0] data_mem_addr[1]
+ data_mem_addr[2] data_mem_addr[3] data_mem_addr[4] data_mem_addr[5] data_mem_addr[6]
+ data_mem_addr[7] hlt instr[0] instr[10] instr[11] instr[12] instr[13] instr[14]
+ instr[15] instr[1] instr[2] instr[3] instr[4] instr[5] instr[6] instr[7] instr[8]
+ instr[9] instr_mem_addr[0] instr_mem_addr[10] instr_mem_addr[11] instr_mem_addr[12]
+ instr_mem_addr[1] instr_mem_addr[2] instr_mem_addr[3] instr_mem_addr[4] instr_mem_addr[5]
+ instr_mem_addr[6] instr_mem_addr[7] instr_mem_addr[8] instr_mem_addr[9] read_data[0]
+ read_data[10] read_data[11] read_data[12] read_data[13] read_data[14] read_data[15]
+ read_data[1] read_data[2] read_data[3] read_data[4] read_data[5] read_data[6] read_data[7]
+ read_data[8] read_data[9] reset start vccd1 vssd1 write_data[0] write_data[10] write_data[11]
+ write_data[12] write_data[13] write_data[14] write_data[15] write_data[1] write_data[2]
+ write_data[3] write_data[4] write_data[5] write_data[6] write_data[7] write_data[8]
+ write_data[9]
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xinstr_memory4 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory4/addr1[0] instr_memory4/addr1[1] instr_memory4/addr1[2]
+ instr_memory4/addr1[3] instr_memory4/addr1[4] instr_memory4/addr1[5] instr_memory4/addr1[6]
+ instr_memory4/addr1[7] instr_memory4/addr1[8] instr_mem_csb\[4\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data4\[0\]
+ instr_read_data4\[1\] instr_read_data4\[2\] instr_read_data4\[3\] instr_read_data4\[4\]
+ instr_read_data4\[5\] instr_read_data4\[6\] instr_read_data4\[7\] instr_read_data4\[8\]
+ instr_read_data4\[9\] instr_read_data4\[10\] instr_read_data4\[11\] instr_read_data4\[12\]
+ instr_read_data4\[13\] instr_read_data4\[14\] instr_read_data4\[15\] instr_read_data4\[16\]
+ instr_read_data4\[17\] instr_read_data4\[18\] instr_read_data4\[19\] instr_read_data4\[20\]
+ instr_read_data4\[21\] instr_read_data4\[22\] instr_read_data4\[23\] instr_read_data4\[24\]
+ instr_read_data4\[25\] instr_read_data4\[26\] instr_read_data4\[27\] instr_read_data4\[28\]
+ instr_read_data4\[29\] instr_read_data4\[30\] instr_read_data4\[31\] instr_memory4/dout1[0]
+ instr_memory4/dout1[1] instr_memory4/dout1[2] instr_memory4/dout1[3] instr_memory4/dout1[4]
+ instr_memory4/dout1[5] instr_memory4/dout1[6] instr_memory4/dout1[7] instr_memory4/dout1[8]
+ instr_memory4/dout1[9] instr_memory4/dout1[10] instr_memory4/dout1[11] instr_memory4/dout1[12]
+ instr_memory4/dout1[13] instr_memory4/dout1[14] instr_memory4/dout1[15] instr_memory4/dout1[16]
+ instr_memory4/dout1[17] instr_memory4/dout1[18] instr_memory4/dout1[19] instr_memory4/dout1[20]
+ instr_memory4/dout1[21] instr_memory4/dout1[22] instr_memory4/dout1[23] instr_memory4/dout1[24]
+ instr_memory4/dout1[25] instr_memory4/dout1[26] instr_memory4/dout1[27] instr_memory4/dout1[28]
+ instr_memory4/dout1[29] instr_memory4/dout1[30] instr_memory4/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
Xinstr_memory5 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory5/addr1[0] instr_memory5/addr1[1] instr_memory5/addr1[2]
+ instr_memory5/addr1[3] instr_memory5/addr1[4] instr_memory5/addr1[5] instr_memory5/addr1[6]
+ instr_memory5/addr1[7] instr_memory5/addr1[8] instr_mem_csb\[5\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data5\[0\]
+ instr_read_data5\[1\] instr_read_data5\[2\] instr_read_data5\[3\] instr_read_data5\[4\]
+ instr_read_data5\[5\] instr_read_data5\[6\] instr_read_data5\[7\] instr_read_data5\[8\]
+ instr_read_data5\[9\] instr_read_data5\[10\] instr_read_data5\[11\] instr_read_data5\[12\]
+ instr_read_data5\[13\] instr_read_data5\[14\] instr_read_data5\[15\] instr_read_data5\[16\]
+ instr_read_data5\[17\] instr_read_data5\[18\] instr_read_data5\[19\] instr_read_data5\[20\]
+ instr_read_data5\[21\] instr_read_data5\[22\] instr_read_data5\[23\] instr_read_data5\[24\]
+ instr_read_data5\[25\] instr_read_data5\[26\] instr_read_data5\[27\] instr_read_data5\[28\]
+ instr_read_data5\[29\] instr_read_data5\[30\] instr_read_data5\[31\] instr_memory5/dout1[0]
+ instr_memory5/dout1[1] instr_memory5/dout1[2] instr_memory5/dout1[3] instr_memory5/dout1[4]
+ instr_memory5/dout1[5] instr_memory5/dout1[6] instr_memory5/dout1[7] instr_memory5/dout1[8]
+ instr_memory5/dout1[9] instr_memory5/dout1[10] instr_memory5/dout1[11] instr_memory5/dout1[12]
+ instr_memory5/dout1[13] instr_memory5/dout1[14] instr_memory5/dout1[15] instr_memory5/dout1[16]
+ instr_memory5/dout1[17] instr_memory5/dout1[18] instr_memory5/dout1[19] instr_memory5/dout1[20]
+ instr_memory5/dout1[21] instr_memory5/dout1[22] instr_memory5/dout1[23] instr_memory5/dout1[24]
+ instr_memory5/dout1[25] instr_memory5/dout1[26] instr_memory5/dout1[27] instr_memory5/dout1[28]
+ instr_memory5/dout1[29] instr_memory5/dout1[30] instr_memory5/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
Xinstr_memory6 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory6/addr1[0] instr_memory6/addr1[1] instr_memory6/addr1[2]
+ instr_memory6/addr1[3] instr_memory6/addr1[4] instr_memory6/addr1[5] instr_memory6/addr1[6]
+ instr_memory6/addr1[7] instr_memory6/addr1[8] instr_mem_csb\[6\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data6\[0\]
+ instr_read_data6\[1\] instr_read_data6\[2\] instr_read_data6\[3\] instr_read_data6\[4\]
+ instr_read_data6\[5\] instr_read_data6\[6\] instr_read_data6\[7\] instr_read_data6\[8\]
+ instr_read_data6\[9\] instr_read_data6\[10\] instr_read_data6\[11\] instr_read_data6\[12\]
+ instr_read_data6\[13\] instr_read_data6\[14\] instr_read_data6\[15\] instr_read_data6\[16\]
+ instr_read_data6\[17\] instr_read_data6\[18\] instr_read_data6\[19\] instr_read_data6\[20\]
+ instr_read_data6\[21\] instr_read_data6\[22\] instr_read_data6\[23\] instr_read_data6\[24\]
+ instr_read_data6\[25\] instr_read_data6\[26\] instr_read_data6\[27\] instr_read_data6\[28\]
+ instr_read_data6\[29\] instr_read_data6\[30\] instr_read_data6\[31\] instr_memory6/dout1[0]
+ instr_memory6/dout1[1] instr_memory6/dout1[2] instr_memory6/dout1[3] instr_memory6/dout1[4]
+ instr_memory6/dout1[5] instr_memory6/dout1[6] instr_memory6/dout1[7] instr_memory6/dout1[8]
+ instr_memory6/dout1[9] instr_memory6/dout1[10] instr_memory6/dout1[11] instr_memory6/dout1[12]
+ instr_memory6/dout1[13] instr_memory6/dout1[14] instr_memory6/dout1[15] instr_memory6/dout1[16]
+ instr_memory6/dout1[17] instr_memory6/dout1[18] instr_memory6/dout1[19] instr_memory6/dout1[20]
+ instr_memory6/dout1[21] instr_memory6/dout1[22] instr_memory6/dout1[23] instr_memory6/dout1[24]
+ instr_memory6/dout1[25] instr_memory6/dout1[26] instr_memory6/dout1[27] instr_memory6/dout1[28]
+ instr_memory6/dout1[29] instr_memory6/dout1[30] instr_memory6/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
Xdata_memory data_write_data\[0\] data_write_data\[1\] data_write_data\[2\] data_write_data\[3\]
+ data_write_data\[4\] data_write_data\[5\] data_write_data\[6\] data_write_data\[7\]
+ data_write_data\[8\] data_write_data\[9\] data_write_data\[10\] data_write_data\[11\]
+ data_write_data\[12\] data_write_data\[13\] data_write_data\[14\] data_write_data\[15\]
+ data_memory/din0[16] data_memory/din0[17] data_memory/din0[18] data_memory/din0[19]
+ data_memory/din0[20] data_memory/din0[21] data_memory/din0[22] data_memory/din0[23]
+ data_memory/din0[24] data_memory/din0[25] data_memory/din0[26] data_memory/din0[27]
+ data_memory/din0[28] data_memory/din0[29] data_memory/din0[30] data_memory/din0[31]
+ data_mem_addr\[0\] data_mem_addr\[1\] data_mem_addr\[2\] data_mem_addr\[3\] data_mem_addr\[4\]
+ data_mem_addr\[5\] data_mem_addr\[6\] data_mem_addr\[7\] low data_memory/addr1[0]
+ data_memory/addr1[1] data_memory/addr1[2] data_memory/addr1[3] data_memory/addr1[4]
+ data_memory/addr1[5] data_memory/addr1[6] data_memory/addr1[7] data_memory/addr1[8]
+ data_mem_csb low dataw_enb clk clk data_wmask\[0\] data_wmask\[1\] data_wmask\[2\]
+ data_wmask\[3\] data_read_data\[0\] data_read_data\[1\] data_read_data\[2\] data_read_data\[3\]
+ data_read_data\[4\] data_read_data\[5\] data_read_data\[6\] data_read_data\[7\]
+ data_read_data\[8\] data_read_data\[9\] data_read_data\[10\] data_read_data\[11\]
+ data_read_data\[12\] data_read_data\[13\] data_read_data\[14\] data_read_data\[15\]
+ data_memory/dout0[16] data_memory/dout0[17] data_memory/dout0[18] data_memory/dout0[19]
+ data_memory/dout0[20] data_memory/dout0[21] data_memory/dout0[22] data_memory/dout0[23]
+ data_memory/dout0[24] data_memory/dout0[25] data_memory/dout0[26] data_memory/dout0[27]
+ data_memory/dout0[28] data_memory/dout0[29] data_memory/dout0[30] data_memory/dout0[31]
+ data_memory/dout1[0] data_memory/dout1[1] data_memory/dout1[2] data_memory/dout1[3]
+ data_memory/dout1[4] data_memory/dout1[5] data_memory/dout1[6] data_memory/dout1[7]
+ data_memory/dout1[8] data_memory/dout1[9] data_memory/dout1[10] data_memory/dout1[11]
+ data_memory/dout1[12] data_memory/dout1[13] data_memory/dout1[14] data_memory/dout1[15]
+ data_memory/dout1[16] data_memory/dout1[17] data_memory/dout1[18] data_memory/dout1[19]
+ data_memory/dout1[20] data_memory/dout1[21] data_memory/dout1[22] data_memory/dout1[23]
+ data_memory/dout1[24] data_memory/dout1[25] data_memory/dout1[26] data_memory/dout1[27]
+ data_memory/dout1[28] data_memory/dout1[29] data_memory/dout1[30] data_memory/dout1[31]
+ vccd1 vssd1 sky130_sram_2kbyte_1rw1r_32x512_8
Xinstr_memory7 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory7/addr1[0] instr_memory7/addr1[1] instr_memory7/addr1[2]
+ instr_memory7/addr1[3] instr_memory7/addr1[4] instr_memory7/addr1[5] instr_memory7/addr1[6]
+ instr_memory7/addr1[7] instr_memory7/addr1[8] instr_mem_csb\[7\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data7\[0\]
+ instr_read_data7\[1\] instr_read_data7\[2\] instr_read_data7\[3\] instr_read_data7\[4\]
+ instr_read_data7\[5\] instr_read_data7\[6\] instr_read_data7\[7\] instr_read_data7\[8\]
+ instr_read_data7\[9\] instr_read_data7\[10\] instr_read_data7\[11\] instr_read_data7\[12\]
+ instr_read_data7\[13\] instr_read_data7\[14\] instr_read_data7\[15\] instr_read_data7\[16\]
+ instr_read_data7\[17\] instr_read_data7\[18\] instr_read_data7\[19\] instr_read_data7\[20\]
+ instr_read_data7\[21\] instr_read_data7\[22\] instr_read_data7\[23\] instr_read_data7\[24\]
+ instr_read_data7\[25\] instr_read_data7\[26\] instr_read_data7\[27\] instr_read_data7\[28\]
+ instr_read_data7\[29\] instr_read_data7\[30\] instr_read_data7\[31\] instr_memory7/dout1[0]
+ instr_memory7/dout1[1] instr_memory7/dout1[2] instr_memory7/dout1[3] instr_memory7/dout1[4]
+ instr_memory7/dout1[5] instr_memory7/dout1[6] instr_memory7/dout1[7] instr_memory7/dout1[8]
+ instr_memory7/dout1[9] instr_memory7/dout1[10] instr_memory7/dout1[11] instr_memory7/dout1[12]
+ instr_memory7/dout1[13] instr_memory7/dout1[14] instr_memory7/dout1[15] instr_memory7/dout1[16]
+ instr_memory7/dout1[17] instr_memory7/dout1[18] instr_memory7/dout1[19] instr_memory7/dout1[20]
+ instr_memory7/dout1[21] instr_memory7/dout1[22] instr_memory7/dout1[23] instr_memory7/dout1[24]
+ instr_memory7/dout1[25] instr_memory7/dout1[26] instr_memory7/dout1[27] instr_memory7/dout1[28]
+ instr_memory7/dout1[29] instr_memory7/dout1[30] instr_memory7/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
XIO_interface Serial_input Serial_output clk data_mem_addr\[0\] data_mem_addr\[1\]
+ data_mem_addr\[2\] data_mem_addr\[3\] data_mem_addr\[4\] data_mem_addr\[5\] data_mem_addr\[6\]
+ data_mem_addr\[7\] data_mem_csb data_read_data\[0\] data_read_data\[10\] data_read_data\[11\]
+ data_read_data\[12\] data_read_data\[13\] data_read_data\[14\] data_read_data\[15\]
+ data_read_data\[1\] data_read_data\[2\] data_read_data\[3\] data_read_data\[4\]
+ data_read_data\[5\] data_read_data\[6\] data_read_data\[7\] data_read_data\[8\]
+ data_read_data\[9\] data_wmask\[0\] data_wmask\[1\] data_wmask\[2\] data_wmask\[3\]
+ data_write_data\[0\] data_write_data\[10\] data_write_data\[11\] data_write_data\[12\]
+ data_write_data\[13\] data_write_data\[14\] data_write_data\[15\] data_write_data\[1\]
+ data_write_data\[2\] data_write_data\[3\] data_write_data\[4\] data_write_data\[5\]
+ data_write_data\[6\] data_write_data\[7\] data_write_data\[8\] data_write_data\[9\]
+ dataw_enb IO_interface/high hlt instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\]
+ instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\] instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\]
+ instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\] instr_mem_addr_9bit\[8\] instr_mem_csb\[7\]
+ instr_mem_csb\[6\] instr_mem_csb\[5\] instr_mem_csb\[4\] instr_mem_csb\[3\] instr_mem_csb\[2\]
+ instr_mem_csb\[1\] instr_mem_csb\[0\] instr_read_data0\[0\] instr_read_data0\[10\]
+ instr_read_data0\[11\] instr_read_data0\[12\] instr_read_data0\[13\] instr_read_data0\[14\]
+ instr_read_data0\[15\] instr_read_data0\[16\] instr_read_data0\[17\] instr_read_data0\[18\]
+ instr_read_data0\[19\] instr_read_data0\[1\] instr_read_data0\[20\] instr_read_data0\[21\]
+ instr_read_data0\[22\] instr_read_data0\[23\] instr_read_data0\[24\] instr_read_data0\[25\]
+ instr_read_data0\[26\] instr_read_data0\[27\] instr_read_data0\[28\] instr_read_data0\[29\]
+ instr_read_data0\[2\] instr_read_data0\[30\] instr_read_data0\[31\] instr_read_data0\[3\]
+ instr_read_data0\[4\] instr_read_data0\[5\] instr_read_data0\[6\] instr_read_data0\[7\]
+ instr_read_data0\[8\] instr_read_data0\[9\] instr_read_data1\[0\] instr_read_data1\[10\]
+ instr_read_data1\[11\] instr_read_data1\[12\] instr_read_data1\[13\] instr_read_data1\[14\]
+ instr_read_data1\[15\] instr_read_data1\[16\] instr_read_data1\[17\] instr_read_data1\[18\]
+ instr_read_data1\[19\] instr_read_data1\[1\] instr_read_data1\[20\] instr_read_data1\[21\]
+ instr_read_data1\[22\] instr_read_data1\[23\] instr_read_data1\[24\] instr_read_data1\[25\]
+ instr_read_data1\[26\] instr_read_data1\[27\] instr_read_data1\[28\] instr_read_data1\[29\]
+ instr_read_data1\[2\] instr_read_data1\[30\] instr_read_data1\[31\] instr_read_data1\[3\]
+ instr_read_data1\[4\] instr_read_data1\[5\] instr_read_data1\[6\] instr_read_data1\[7\]
+ instr_read_data1\[8\] instr_read_data1\[9\] instr_read_data2\[0\] instr_read_data2\[10\]
+ instr_read_data2\[11\] instr_read_data2\[12\] instr_read_data2\[13\] instr_read_data2\[14\]
+ instr_read_data2\[15\] instr_read_data2\[16\] instr_read_data2\[17\] instr_read_data2\[18\]
+ instr_read_data2\[19\] instr_read_data2\[1\] instr_read_data2\[20\] instr_read_data2\[21\]
+ instr_read_data2\[22\] instr_read_data2\[23\] instr_read_data2\[24\] instr_read_data2\[25\]
+ instr_read_data2\[26\] instr_read_data2\[27\] instr_read_data2\[28\] instr_read_data2\[29\]
+ instr_read_data2\[2\] instr_read_data2\[30\] instr_read_data2\[31\] instr_read_data2\[3\]
+ instr_read_data2\[4\] instr_read_data2\[5\] instr_read_data2\[6\] instr_read_data2\[7\]
+ instr_read_data2\[8\] instr_read_data2\[9\] instr_read_data3\[0\] instr_read_data3\[10\]
+ instr_read_data3\[11\] instr_read_data3\[12\] instr_read_data3\[13\] instr_read_data3\[14\]
+ instr_read_data3\[15\] instr_read_data3\[16\] instr_read_data3\[17\] instr_read_data3\[18\]
+ instr_read_data3\[19\] instr_read_data3\[1\] instr_read_data3\[20\] instr_read_data3\[21\]
+ instr_read_data3\[22\] instr_read_data3\[23\] instr_read_data3\[24\] instr_read_data3\[25\]
+ instr_read_data3\[26\] instr_read_data3\[27\] instr_read_data3\[28\] instr_read_data3\[29\]
+ instr_read_data3\[2\] instr_read_data3\[30\] instr_read_data3\[31\] instr_read_data3\[3\]
+ instr_read_data3\[4\] instr_read_data3\[5\] instr_read_data3\[6\] instr_read_data3\[7\]
+ instr_read_data3\[8\] instr_read_data3\[9\] instr_read_data4\[0\] instr_read_data4\[10\]
+ instr_read_data4\[11\] instr_read_data4\[12\] instr_read_data4\[13\] instr_read_data4\[14\]
+ instr_read_data4\[15\] instr_read_data4\[16\] instr_read_data4\[17\] instr_read_data4\[18\]
+ instr_read_data4\[19\] instr_read_data4\[1\] instr_read_data4\[20\] instr_read_data4\[21\]
+ instr_read_data4\[22\] instr_read_data4\[23\] instr_read_data4\[24\] instr_read_data4\[25\]
+ instr_read_data4\[26\] instr_read_data4\[27\] instr_read_data4\[28\] instr_read_data4\[29\]
+ instr_read_data4\[2\] instr_read_data4\[30\] instr_read_data4\[31\] instr_read_data4\[3\]
+ instr_read_data4\[4\] instr_read_data4\[5\] instr_read_data4\[6\] instr_read_data4\[7\]
+ instr_read_data4\[8\] instr_read_data4\[9\] instr_read_data5\[0\] instr_read_data5\[10\]
+ instr_read_data5\[11\] instr_read_data5\[12\] instr_read_data5\[13\] instr_read_data5\[14\]
+ instr_read_data5\[15\] instr_read_data5\[16\] instr_read_data5\[17\] instr_read_data5\[18\]
+ instr_read_data5\[19\] instr_read_data5\[1\] instr_read_data5\[20\] instr_read_data5\[21\]
+ instr_read_data5\[22\] instr_read_data5\[23\] instr_read_data5\[24\] instr_read_data5\[25\]
+ instr_read_data5\[26\] instr_read_data5\[27\] instr_read_data5\[28\] instr_read_data5\[29\]
+ instr_read_data5\[2\] instr_read_data5\[30\] instr_read_data5\[31\] instr_read_data5\[3\]
+ instr_read_data5\[4\] instr_read_data5\[5\] instr_read_data5\[6\] instr_read_data5\[7\]
+ instr_read_data5\[8\] instr_read_data5\[9\] instr_read_data6\[0\] instr_read_data6\[10\]
+ instr_read_data6\[11\] instr_read_data6\[12\] instr_read_data6\[13\] instr_read_data6\[14\]
+ instr_read_data6\[15\] instr_read_data6\[16\] instr_read_data6\[17\] instr_read_data6\[18\]
+ instr_read_data6\[19\] instr_read_data6\[1\] instr_read_data6\[20\] instr_read_data6\[21\]
+ instr_read_data6\[22\] instr_read_data6\[23\] instr_read_data6\[24\] instr_read_data6\[25\]
+ instr_read_data6\[26\] instr_read_data6\[27\] instr_read_data6\[28\] instr_read_data6\[29\]
+ instr_read_data6\[2\] instr_read_data6\[30\] instr_read_data6\[31\] instr_read_data6\[3\]
+ instr_read_data6\[4\] instr_read_data6\[5\] instr_read_data6\[6\] instr_read_data6\[7\]
+ instr_read_data6\[8\] instr_read_data6\[9\] instr_read_data7\[0\] instr_read_data7\[10\]
+ instr_read_data7\[11\] instr_read_data7\[12\] instr_read_data7\[13\] instr_read_data7\[14\]
+ instr_read_data7\[15\] instr_read_data7\[16\] instr_read_data7\[17\] instr_read_data7\[18\]
+ instr_read_data7\[19\] instr_read_data7\[1\] instr_read_data7\[20\] instr_read_data7\[21\]
+ instr_read_data7\[22\] instr_read_data7\[23\] instr_read_data7\[24\] instr_read_data7\[25\]
+ instr_read_data7\[26\] instr_read_data7\[27\] instr_read_data7\[28\] instr_read_data7\[29\]
+ instr_read_data7\[2\] instr_read_data7\[30\] instr_read_data7\[31\] instr_read_data7\[3\]
+ instr_read_data7\[4\] instr_read_data7\[5\] instr_read_data7\[6\] instr_read_data7\[7\]
+ instr_read_data7\[8\] instr_read_data7\[9\] instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\]
+ instr_wmask\[3\] instr_write_data\[0\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\] instr_write_data\[4\]
+ instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\] instr_write_data\[8\]
+ instr_write_data\[9\] instrw_enb io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] user_irq[0] user_irq[1] user_irq[2] la_data_in[0] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] low reset
+ start uP_data_mem_addr\[0\] uP_data_mem_addr\[1\] uP_data_mem_addr\[2\] uP_data_mem_addr\[3\]
+ uP_data_mem_addr\[4\] uP_data_mem_addr\[5\] uP_data_mem_addr\[6\] uP_data_mem_addr\[7\]
+ uP_dataw_en uP_instr\[0\] uP_instr\[10\] uP_instr\[11\] uP_instr\[12\] uP_instr\[13\]
+ uP_instr\[14\] uP_instr\[15\] uP_instr\[1\] uP_instr\[2\] uP_instr\[3\] uP_instr\[4\]
+ uP_instr\[5\] uP_instr\[6\] uP_instr\[7\] uP_instr\[8\] uP_instr\[9\] uP_instr_mem_addr\[0\]
+ uP_instr_mem_addr\[10\] uP_instr_mem_addr\[11\] uP_instr_mem_addr\[12\] uP_instr_mem_addr\[1\]
+ uP_instr_mem_addr\[2\] uP_instr_mem_addr\[3\] uP_instr_mem_addr\[4\] uP_instr_mem_addr\[5\]
+ uP_instr_mem_addr\[6\] uP_instr_mem_addr\[7\] uP_instr_mem_addr\[8\] uP_instr_mem_addr\[9\]
+ uP_read_data\[0\] uP_read_data\[10\] uP_read_data\[11\] uP_read_data\[12\] uP_read_data\[13\]
+ uP_read_data\[14\] uP_read_data\[15\] uP_read_data\[1\] uP_read_data\[2\] uP_read_data\[3\]
+ uP_read_data\[4\] uP_read_data\[5\] uP_read_data\[6\] uP_read_data\[7\] uP_read_data\[8\]
+ uP_read_data\[9\] uP_write_data\[0\] uP_write_data\[10\] uP_write_data\[11\] uP_write_data\[12\]
+ uP_write_data\[13\] uP_write_data\[14\] uP_write_data\[15\] uP_write_data\[1\] uP_write_data\[2\]
+ uP_write_data\[3\] uP_write_data\[4\] uP_write_data\[5\] uP_write_data\[6\] uP_write_data\[7\]
+ uP_write_data\[8\] uP_write_data\[9\] vccd1 vssd1 wb_clk_i wb_rst_i io_interface
Xinstr_memory0 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory0/addr1[0] instr_memory0/addr1[1] instr_memory0/addr1[2]
+ instr_memory0/addr1[3] instr_memory0/addr1[4] instr_memory0/addr1[5] instr_memory0/addr1[6]
+ instr_memory0/addr1[7] instr_memory0/addr1[8] instr_mem_csb\[0\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data0\[0\]
+ instr_read_data0\[1\] instr_read_data0\[2\] instr_read_data0\[3\] instr_read_data0\[4\]
+ instr_read_data0\[5\] instr_read_data0\[6\] instr_read_data0\[7\] instr_read_data0\[8\]
+ instr_read_data0\[9\] instr_read_data0\[10\] instr_read_data0\[11\] instr_read_data0\[12\]
+ instr_read_data0\[13\] instr_read_data0\[14\] instr_read_data0\[15\] instr_read_data0\[16\]
+ instr_read_data0\[17\] instr_read_data0\[18\] instr_read_data0\[19\] instr_read_data0\[20\]
+ instr_read_data0\[21\] instr_read_data0\[22\] instr_read_data0\[23\] instr_read_data0\[24\]
+ instr_read_data0\[25\] instr_read_data0\[26\] instr_read_data0\[27\] instr_read_data0\[28\]
+ instr_read_data0\[29\] instr_read_data0\[30\] instr_read_data0\[31\] instr_memory0/dout1[0]
+ instr_memory0/dout1[1] instr_memory0/dout1[2] instr_memory0/dout1[3] instr_memory0/dout1[4]
+ instr_memory0/dout1[5] instr_memory0/dout1[6] instr_memory0/dout1[7] instr_memory0/dout1[8]
+ instr_memory0/dout1[9] instr_memory0/dout1[10] instr_memory0/dout1[11] instr_memory0/dout1[12]
+ instr_memory0/dout1[13] instr_memory0/dout1[14] instr_memory0/dout1[15] instr_memory0/dout1[16]
+ instr_memory0/dout1[17] instr_memory0/dout1[18] instr_memory0/dout1[19] instr_memory0/dout1[20]
+ instr_memory0/dout1[21] instr_memory0/dout1[22] instr_memory0/dout1[23] instr_memory0/dout1[24]
+ instr_memory0/dout1[25] instr_memory0/dout1[26] instr_memory0/dout1[27] instr_memory0/dout1[28]
+ instr_memory0/dout1[29] instr_memory0/dout1[30] instr_memory0/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
Xinstr_memory1 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory1/addr1[0] instr_memory1/addr1[1] instr_memory1/addr1[2]
+ instr_memory1/addr1[3] instr_memory1/addr1[4] instr_memory1/addr1[5] instr_memory1/addr1[6]
+ instr_memory1/addr1[7] instr_memory1/addr1[8] instr_mem_csb\[1\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data1\[0\]
+ instr_read_data1\[1\] instr_read_data1\[2\] instr_read_data1\[3\] instr_read_data1\[4\]
+ instr_read_data1\[5\] instr_read_data1\[6\] instr_read_data1\[7\] instr_read_data1\[8\]
+ instr_read_data1\[9\] instr_read_data1\[10\] instr_read_data1\[11\] instr_read_data1\[12\]
+ instr_read_data1\[13\] instr_read_data1\[14\] instr_read_data1\[15\] instr_read_data1\[16\]
+ instr_read_data1\[17\] instr_read_data1\[18\] instr_read_data1\[19\] instr_read_data1\[20\]
+ instr_read_data1\[21\] instr_read_data1\[22\] instr_read_data1\[23\] instr_read_data1\[24\]
+ instr_read_data1\[25\] instr_read_data1\[26\] instr_read_data1\[27\] instr_read_data1\[28\]
+ instr_read_data1\[29\] instr_read_data1\[30\] instr_read_data1\[31\] instr_memory1/dout1[0]
+ instr_memory1/dout1[1] instr_memory1/dout1[2] instr_memory1/dout1[3] instr_memory1/dout1[4]
+ instr_memory1/dout1[5] instr_memory1/dout1[6] instr_memory1/dout1[7] instr_memory1/dout1[8]
+ instr_memory1/dout1[9] instr_memory1/dout1[10] instr_memory1/dout1[11] instr_memory1/dout1[12]
+ instr_memory1/dout1[13] instr_memory1/dout1[14] instr_memory1/dout1[15] instr_memory1/dout1[16]
+ instr_memory1/dout1[17] instr_memory1/dout1[18] instr_memory1/dout1[19] instr_memory1/dout1[20]
+ instr_memory1/dout1[21] instr_memory1/dout1[22] instr_memory1/dout1[23] instr_memory1/dout1[24]
+ instr_memory1/dout1[25] instr_memory1/dout1[26] instr_memory1/dout1[27] instr_memory1/dout1[28]
+ instr_memory1/dout1[29] instr_memory1/dout1[30] instr_memory1/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
Xinstr_memory2 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory2/addr1[0] instr_memory2/addr1[1] instr_memory2/addr1[2]
+ instr_memory2/addr1[3] instr_memory2/addr1[4] instr_memory2/addr1[5] instr_memory2/addr1[6]
+ instr_memory2/addr1[7] instr_memory2/addr1[8] instr_mem_csb\[2\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data2\[0\]
+ instr_read_data2\[1\] instr_read_data2\[2\] instr_read_data2\[3\] instr_read_data2\[4\]
+ instr_read_data2\[5\] instr_read_data2\[6\] instr_read_data2\[7\] instr_read_data2\[8\]
+ instr_read_data2\[9\] instr_read_data2\[10\] instr_read_data2\[11\] instr_read_data2\[12\]
+ instr_read_data2\[13\] instr_read_data2\[14\] instr_read_data2\[15\] instr_read_data2\[16\]
+ instr_read_data2\[17\] instr_read_data2\[18\] instr_read_data2\[19\] instr_read_data2\[20\]
+ instr_read_data2\[21\] instr_read_data2\[22\] instr_read_data2\[23\] instr_read_data2\[24\]
+ instr_read_data2\[25\] instr_read_data2\[26\] instr_read_data2\[27\] instr_read_data2\[28\]
+ instr_read_data2\[29\] instr_read_data2\[30\] instr_read_data2\[31\] instr_memory2/dout1[0]
+ instr_memory2/dout1[1] instr_memory2/dout1[2] instr_memory2/dout1[3] instr_memory2/dout1[4]
+ instr_memory2/dout1[5] instr_memory2/dout1[6] instr_memory2/dout1[7] instr_memory2/dout1[8]
+ instr_memory2/dout1[9] instr_memory2/dout1[10] instr_memory2/dout1[11] instr_memory2/dout1[12]
+ instr_memory2/dout1[13] instr_memory2/dout1[14] instr_memory2/dout1[15] instr_memory2/dout1[16]
+ instr_memory2/dout1[17] instr_memory2/dout1[18] instr_memory2/dout1[19] instr_memory2/dout1[20]
+ instr_memory2/dout1[21] instr_memory2/dout1[22] instr_memory2/dout1[23] instr_memory2/dout1[24]
+ instr_memory2/dout1[25] instr_memory2/dout1[26] instr_memory2/dout1[27] instr_memory2/dout1[28]
+ instr_memory2/dout1[29] instr_memory2/dout1[30] instr_memory2/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
XuP uP_dataw_en Serial_input Serial_output clk uP_data_mem_addr\[0\] uP_data_mem_addr\[1\]
+ uP_data_mem_addr\[2\] uP_data_mem_addr\[3\] uP_data_mem_addr\[4\] uP_data_mem_addr\[5\]
+ uP_data_mem_addr\[6\] uP_data_mem_addr\[7\] hlt uP_instr\[0\] uP_instr\[10\] uP_instr\[11\]
+ uP_instr\[12\] uP_instr\[13\] uP_instr\[14\] uP_instr\[15\] uP_instr\[1\] uP_instr\[2\]
+ uP_instr\[3\] uP_instr\[4\] uP_instr\[5\] uP_instr\[6\] uP_instr\[7\] uP_instr\[8\]
+ uP_instr\[9\] uP_instr_mem_addr\[0\] uP_instr_mem_addr\[10\] uP_instr_mem_addr\[11\]
+ uP_instr_mem_addr\[12\] uP_instr_mem_addr\[1\] uP_instr_mem_addr\[2\] uP_instr_mem_addr\[3\]
+ uP_instr_mem_addr\[4\] uP_instr_mem_addr\[5\] uP_instr_mem_addr\[6\] uP_instr_mem_addr\[7\]
+ uP_instr_mem_addr\[8\] uP_instr_mem_addr\[9\] uP_read_data\[0\] uP_read_data\[10\]
+ uP_read_data\[11\] uP_read_data\[12\] uP_read_data\[13\] uP_read_data\[14\] uP_read_data\[15\]
+ uP_read_data\[1\] uP_read_data\[2\] uP_read_data\[3\] uP_read_data\[4\] uP_read_data\[5\]
+ uP_read_data\[6\] uP_read_data\[7\] uP_read_data\[8\] uP_read_data\[9\] reset start
+ vccd1 vssd1 uP_write_data\[0\] uP_write_data\[10\] uP_write_data\[11\] uP_write_data\[12\]
+ uP_write_data\[13\] uP_write_data\[14\] uP_write_data\[15\] uP_write_data\[1\] uP_write_data\[2\]
+ uP_write_data\[3\] uP_write_data\[4\] uP_write_data\[5\] uP_write_data\[6\] uP_write_data\[7\]
+ uP_write_data\[8\] uP_write_data\[9\] processor
Xinstr_memory3 instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_write_data\[0\] instr_write_data\[1\] instr_write_data\[2\] instr_write_data\[3\]
+ instr_write_data\[4\] instr_write_data\[5\] instr_write_data\[6\] instr_write_data\[7\]
+ instr_write_data\[8\] instr_write_data\[9\] instr_write_data\[10\] instr_write_data\[11\]
+ instr_write_data\[12\] instr_write_data\[13\] instr_write_data\[14\] instr_write_data\[15\]
+ instr_mem_addr_9bit\[0\] instr_mem_addr_9bit\[1\] instr_mem_addr_9bit\[2\] instr_mem_addr_9bit\[3\]
+ instr_mem_addr_9bit\[4\] instr_mem_addr_9bit\[5\] instr_mem_addr_9bit\[6\] instr_mem_addr_9bit\[7\]
+ instr_mem_addr_9bit\[8\] instr_memory3/addr1[0] instr_memory3/addr1[1] instr_memory3/addr1[2]
+ instr_memory3/addr1[3] instr_memory3/addr1[4] instr_memory3/addr1[5] instr_memory3/addr1[6]
+ instr_memory3/addr1[7] instr_memory3/addr1[8] instr_mem_csb\[3\] low instrw_enb
+ clk clk instr_wmask\[0\] instr_wmask\[1\] instr_wmask\[2\] instr_wmask\[3\] instr_read_data3\[0\]
+ instr_read_data3\[1\] instr_read_data3\[2\] instr_read_data3\[3\] instr_read_data3\[4\]
+ instr_read_data3\[5\] instr_read_data3\[6\] instr_read_data3\[7\] instr_read_data3\[8\]
+ instr_read_data3\[9\] instr_read_data3\[10\] instr_read_data3\[11\] instr_read_data3\[12\]
+ instr_read_data3\[13\] instr_read_data3\[14\] instr_read_data3\[15\] instr_read_data3\[16\]
+ instr_read_data3\[17\] instr_read_data3\[18\] instr_read_data3\[19\] instr_read_data3\[20\]
+ instr_read_data3\[21\] instr_read_data3\[22\] instr_read_data3\[23\] instr_read_data3\[24\]
+ instr_read_data3\[25\] instr_read_data3\[26\] instr_read_data3\[27\] instr_read_data3\[28\]
+ instr_read_data3\[29\] instr_read_data3\[30\] instr_read_data3\[31\] instr_memory3/dout1[0]
+ instr_memory3/dout1[1] instr_memory3/dout1[2] instr_memory3/dout1[3] instr_memory3/dout1[4]
+ instr_memory3/dout1[5] instr_memory3/dout1[6] instr_memory3/dout1[7] instr_memory3/dout1[8]
+ instr_memory3/dout1[9] instr_memory3/dout1[10] instr_memory3/dout1[11] instr_memory3/dout1[12]
+ instr_memory3/dout1[13] instr_memory3/dout1[14] instr_memory3/dout1[15] instr_memory3/dout1[16]
+ instr_memory3/dout1[17] instr_memory3/dout1[18] instr_memory3/dout1[19] instr_memory3/dout1[20]
+ instr_memory3/dout1[21] instr_memory3/dout1[22] instr_memory3/dout1[23] instr_memory3/dout1[24]
+ instr_memory3/dout1[25] instr_memory3/dout1[26] instr_memory3/dout1[27] instr_memory3/dout1[28]
+ instr_memory3/dout1[29] instr_memory3/dout1[30] instr_memory3/dout1[31] vccd1 vssd1
+ sky130_sram_2kbyte_1rw1r_32x512_8
.ends

