magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< locali >>
rect 6053 5476 6087 5492
rect 6053 5426 6087 5442
<< viali >>
rect 6053 5442 6087 5476
<< metal1 >>
rect 6038 5433 6044 5485
rect 6096 5433 6102 5485
rect 2083 -2950 2089 -2898
rect 2141 -2910 2147 -2898
rect 6038 -2910 6044 -2898
rect 2141 -2938 6044 -2910
rect 2141 -2950 2147 -2938
rect 6038 -2950 6044 -2938
rect 6096 -2950 6102 -2898
<< via1 >>
rect 6044 5476 6096 5485
rect 6044 5442 6053 5476
rect 6053 5442 6087 5476
rect 6087 5442 6096 5476
rect 6044 5433 6096 5442
rect 2089 -2950 2141 -2898
rect 6044 -2950 6096 -2898
<< metal2 >>
rect 6044 5485 6096 5491
rect 6044 5427 6096 5433
rect 6056 -2892 6084 5427
rect 2089 -2898 2141 -2892
rect 2089 -2956 2141 -2950
rect 6044 -2898 6096 -2892
rect 6044 -2956 6096 -2950
rect 2101 -3939 2129 -2956
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_0
timestamp 1666464484
transform 1 0 6041 0 1 5426
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1666464484
transform 1 0 2083 0 1 -2956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1666464484
transform 1 0 6038 0 1 5427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1666464484
transform 1 0 6038 0 1 -2956
box 0 0 1 1
<< properties >>
string FIXED_BBOX 2083 -3939 6102 5492
string GDS_END 7324138
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 7323390
<< end >>
